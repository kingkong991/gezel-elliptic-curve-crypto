library ieee;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
library work;
use work.std_logic_arithext.all;


--datapath entity
entity wrapper_pairing is
   port(
      input:in std_logic_vector(162 downto 0);
      start_in:in std_logic;
      next_in:in std_logic;
      output:out std_logic_vector(162 downto 0);
      ready:out std_logic;
      sig_en_out_Xv:out std_logic;
      sig_en_out_Yv:out std_logic;
      sig_en_out_Xp:out std_logic;
      sig_en_out_Yp:out std_logic;
      sig_en_out_Xfa:out std_logic;
      sig_en_out_Yfa:out std_logic;
      sig_en_out_Ga:out std_logic;
      sig_en_out_Gb:out std_logic;
      sig_en_out_Fa:out std_logic;
      sig_en_out_Fb:out std_logic;
      sig_en_out_Fc:out std_logic;
      sig_en_out_Fd:out std_logic;
      sig_en_out_TmpA:out std_logic;
      sig_en_out_TmpB:out std_logic;
      sig_en_out_ToMALU:out std_logic;
      RST : in std_logic;
      CLK : in std_logic
   );
end wrapper_pairing;


--signal declaration
architecture RTL of wrapper_pairing is
signal reg_Xv:std_logic_vector(162 downto 0);
signal reg_Xv_wire:std_logic_vector(162 downto 0);
signal reg_Yv:std_logic_vector(162 downto 0);
signal reg_Yv_wire:std_logic_vector(162 downto 0);
signal reg_Xp:std_logic_vector(162 downto 0);
signal reg_Xp_wire:std_logic_vector(162 downto 0);
signal reg_Yp:std_logic_vector(162 downto 0);
signal reg_Yp_wire:std_logic_vector(162 downto 0);
signal reg_Xfa:std_logic_vector(162 downto 0);
signal reg_Xfa_wire:std_logic_vector(162 downto 0);
signal reg_Yfa:std_logic_vector(162 downto 0);
signal reg_Yfa_wire:std_logic_vector(162 downto 0);
signal reg_Ga:std_logic_vector(162 downto 0);
signal reg_Ga_wire:std_logic_vector(162 downto 0);
signal reg_Gb:std_logic_vector(162 downto 0);
signal reg_Gb_wire:std_logic_vector(162 downto 0);
signal reg_Fa:std_logic_vector(162 downto 0);
signal reg_Fa_wire:std_logic_vector(162 downto 0);
signal reg_Fb:std_logic_vector(162 downto 0);
signal reg_Fb_wire:std_logic_vector(162 downto 0);
signal reg_Fc:std_logic_vector(162 downto 0);
signal reg_Fc_wire:std_logic_vector(162 downto 0);
signal reg_Fd:std_logic_vector(162 downto 0);
signal reg_Fd_wire:std_logic_vector(162 downto 0);
signal reg_TmpA:std_logic_vector(162 downto 0);
signal reg_TmpA_wire:std_logic_vector(162 downto 0);
signal reg_TmpB:std_logic_vector(162 downto 0);
signal reg_TmpB_wire:std_logic_vector(162 downto 0);
signal reg_ToMALU:std_logic_vector(162 downto 0);
signal reg_ToMALU_wire:std_logic_vector(162 downto 0);
signal reg_MALU_ready:std_logic;
signal reg_MALU_ready_wire:std_logic;
signal reg_counter_miller:std_logic_vector(7 downto 0);
signal reg_counter_miller_wire:std_logic_vector(7 downto 0);
signal reg_counter_misc:std_logic_vector(6 downto 0);
signal reg_counter_misc_wire:std_logic_vector(6 downto 0);
signal reg_add:std_logic;
signal reg_add_wire:std_logic;
signal reg_start:std_logic;
signal reg_start_wire:std_logic;
signal reg_next:std_logic;
signal reg_next_wire:std_logic;
signal reg_ready:std_logic;
signal reg_ready_wire:std_logic;
signal sig_MALU_A:std_logic_vector(162 downto 0);
signal sig_MALU_B:std_logic_vector(162 downto 0);
signal sig_MALU_start:std_logic;
signal sig_MALU_mode:std_logic;
signal sig_MALU_plus_one:std_logic;
signal sig_MALU_result:std_logic_vector(162 downto 0);
signal sig_MALU_ready:std_logic;
signal sig_en_Xv:std_logic;
signal sig_en_Yv:std_logic;
signal sig_en_Xp:std_logic;
signal sig_en_Yp:std_logic;
signal sig_en_Xfa:std_logic;
signal sig_en_Yfa:std_logic;
signal sig_en_Ga:std_logic;
signal sig_en_Gb:std_logic;
signal sig_en_Fa:std_logic;
signal sig_en_Fb:std_logic;
signal sig_en_Fc:std_logic;
signal sig_en_Fd:std_logic;
signal sig_en_TmpA:std_logic;
signal sig_en_TmpB:std_logic;
signal sig_en_ToMALU:std_logic;
signal sig_sel_Xv:std_logic_vector(1 downto 0);
signal sig_sel_Yv:std_logic;
signal sig_sel_Xp:std_logic;
signal sig_sel_Yp:std_logic;
signal sig_sel_Xfa:std_logic;
signal sig_sel_Yfa:std_logic;
signal sig_sel_Ga:std_logic;
signal sig_sel_Gb:std_logic;
signal sig_sel_Fa:std_logic;
signal sig_sel_Fb:std_logic;
signal sig_sel_Fc:std_logic;
signal sig_sel_Fd:std_logic;
signal sig_sel_TmpA:std_logic;
signal sig_sel_TmpB:std_logic;
signal sig_sel_ToMALU:std_logic_vector(1 downto 0);
signal sig_to_Xv:std_logic_vector(162 downto 0);
signal sig_to_Yv:std_logic_vector(162 downto 0);
signal sig_to_Xp:std_logic_vector(162 downto 0);
signal sig_to_Yp:std_logic_vector(162 downto 0);
signal sig_to_Xfa:std_logic_vector(162 downto 0);
signal sig_to_Yfa:std_logic_vector(162 downto 0);
signal sig_to_Ga:std_logic_vector(162 downto 0);
signal sig_to_Gb:std_logic_vector(162 downto 0);
signal sig_to_Fa:std_logic_vector(162 downto 0);
signal sig_to_Fb:std_logic_vector(162 downto 0);
signal sig_to_Fc:std_logic_vector(162 downto 0);
signal sig_to_Fd:std_logic_vector(162 downto 0);
signal sig_to_TmpA:std_logic_vector(162 downto 0);
signal sig_to_TmpB:std_logic_vector(162 downto 0);
signal sig_to_ToMALU:std_logic_vector(162 downto 0);
signal sig_from_Xv:std_logic_vector(162 downto 0);
signal sig_from_Yv:std_logic_vector(162 downto 0);
signal sig_from_Xp:std_logic_vector(162 downto 0);
signal sig_from_Yp:std_logic_vector(162 downto 0);
signal sig_from_Xfa:std_logic_vector(162 downto 0);
signal sig_from_Yfa:std_logic_vector(162 downto 0);
signal sig_from_Ga:std_logic_vector(162 downto 0);
signal sig_from_Gb:std_logic_vector(162 downto 0);
signal sig_from_Fa:std_logic_vector(162 downto 0);
signal sig_from_Fb:std_logic_vector(162 downto 0);
signal sig_from_Fc:std_logic_vector(162 downto 0);
signal sig_from_Fd:std_logic_vector(162 downto 0);
signal sig_from_TmpA:std_logic_vector(162 downto 0);
signal sig_from_TmpB:std_logic_vector(162 downto 0);
signal sig_from_ToMALU:std_logic_vector(162 downto 0);
signal sig_from_ToMALUShift:std_logic_vector(162 downto 0);
signal sig_from_Input:std_logic_vector(162 downto 0);
signal sig_0:std_logic;
signal sig_1:std_logic_vector(162 downto 0);
signal sig_2:std_logic_vector(161 downto 0);
signal sig_3:std_logic;
signal sig_4:std_logic_vector(162 downto 0);
signal sig_6:std_logic;
signal sig_8:std_logic;
signal sig_10:std_logic;
signal sig_11:std_logic_vector(162 downto 0);
signal sig_12:std_logic_vector(162 downto 0);
signal sig_13:std_logic;
signal sig_14:std_logic_vector(162 downto 0);
signal sig_15:std_logic;
signal sig_16:std_logic_vector(162 downto 0);
signal sig_17:std_logic;
signal sig_18:std_logic_vector(162 downto 0);
signal sig_19:std_logic;
signal sig_20:std_logic_vector(162 downto 0);
signal sig_21:std_logic;
signal sig_22:std_logic_vector(162 downto 0);
signal sig_23:std_logic;
signal sig_24:std_logic_vector(162 downto 0);
signal sig_25:std_logic;
signal sig_26:std_logic_vector(162 downto 0);
signal sig_27:std_logic;
signal sig_28:std_logic_vector(162 downto 0);
signal sig_29:std_logic;
signal sig_30:std_logic_vector(162 downto 0);
signal sig_31:std_logic;
signal sig_32:std_logic_vector(162 downto 0);
signal sig_33:std_logic;
signal sig_34:std_logic_vector(162 downto 0);
signal sig_35:std_logic;
signal sig_36:std_logic_vector(162 downto 0);
signal sig_37:std_logic;
signal sig_38:std_logic_vector(162 downto 0);
signal sig_40:std_logic;
signal sig_42:std_logic;
signal sig_43:std_logic_vector(162 downto 0);
signal sig_44:std_logic_vector(162 downto 0);
signal sig_56:std_logic_vector(7 downto 0);
signal sig_57:std_logic_vector(6 downto 0);
signal sig_58:std_logic;
signal sig_59:std_logic;
signal sig_60:std_logic;
signal sig_61:std_logic_vector(6 downto 0);
signal sig_62:std_logic_vector(6 downto 0);
signal sig_64:std_logic;
signal sig_65:std_logic;
signal sig_66:std_logic;
signal sig_67:std_logic_vector(162 downto 0);
signal sig_68:std_logic;
signal sig_69:std_logic;
signal sig_70:std_logic;
signal sig_71:std_logic_vector(162 downto 0);
signal sig_72:std_logic;
signal sig_73:std_logic;
signal sig_74:std_logic;
signal sig_75:std_logic_vector(162 downto 0);
signal ready_int:std_logic;
signal output_int:std_logic_vector(162 downto 0);
signal sig_en_out_Xv_int:std_logic;
signal sig_en_out_Yv_int:std_logic;
signal sig_en_out_Xp_int:std_logic;
signal sig_en_out_Yp_int:std_logic;
signal sig_en_out_Xfa_int:std_logic;
signal sig_en_out_Yfa_int:std_logic;
signal sig_en_out_Ga_int:std_logic;
signal sig_en_out_Gb_int:std_logic;
signal sig_en_out_Fa_int:std_logic;
signal sig_en_out_Fb_int:std_logic;
signal sig_en_out_Fc_int:std_logic;
signal sig_en_out_Fd_int:std_logic;
signal sig_en_out_TmpA_int:std_logic;
signal sig_en_out_TmpB_int:std_logic;
signal sig_en_out_ToMALU_int:std_logic;
signal sig_78:std_logic;
signal sig_79:std_logic;
signal sig_80:std_logic;
signal sig_81:std_logic;
signal sig_82:std_logic;
signal sig_83:std_logic;
signal sig_84:std_logic;
signal sig_85:std_logic;
signal sig_86:std_logic;
signal sig_87:std_logic;
signal sig_88:std_logic;
signal sig_89:std_logic;
signal sig_90:std_logic;
signal sig_91:std_logic;
signal sig_92:std_logic;
signal sig_93:std_logic;
signal sig_94:std_logic;
signal sig_95:std_logic;
signal sig_96:std_logic;
signal sig_97:std_logic;
signal sig_98:std_logic;
signal sig_99:std_logic;
signal sig_100:std_logic;
signal sig_101:std_logic;
signal sig_102:std_logic;
signal sig_103:std_logic;
signal sig_104:std_logic;
signal sig_105:std_logic;
signal sig_106:std_logic;
signal sig_107:std_logic;
signal sig_108:std_logic;
signal sig_109:std_logic;
signal sig_110:std_logic;
signal sig_111:std_logic;
signal sig_112:std_logic;
signal sig_113:std_logic;
signal sig_114:std_logic;
signal sig_115:std_logic;
signal sig_116:std_logic;
signal sig_117:std_logic;
signal sig_118:std_logic;
signal sig_119:std_logic;
signal sig_120:std_logic;
signal sig_121:std_logic;
signal sig_122:std_logic;
signal sig_123:std_logic;
signal sig_124:std_logic;
signal sig_125:std_logic;
signal sig_126:std_logic;
signal sig_127:std_logic;
signal sig_128:std_logic;
signal sig_129:std_logic;
signal sig_130:std_logic;
signal sig_131:std_logic;
signal sig_132:std_logic;
signal sig_133:std_logic;
signal sig_134:std_logic;
signal sig_135:std_logic;
signal sig_136:std_logic;
signal sig_137:std_logic;
signal sig_138:std_logic;
signal sig_139:std_logic;
signal sig_140:std_logic;
signal sig_141:std_logic;
signal sig_142:std_logic;
signal sig_143:std_logic;
signal sig_144:std_logic;
signal sig_145:std_logic;
signal sig_146:std_logic;
signal sig_147:std_logic;
signal sig_148:std_logic;
signal sig_149:std_logic;
signal sig_150:std_logic;
signal sig_151:std_logic;
signal sig_152:std_logic;
signal sig_153:std_logic;
signal sig_154:std_logic;
signal sig_155:std_logic;
signal sig_156:std_logic;
signal sig_157:std_logic;
signal sig_158:std_logic;
signal sig_159:std_logic;
signal sig_160:std_logic;
signal sig_161:std_logic;
signal sig_162:std_logic;
signal sig_163:std_logic;
signal sig_164:std_logic;
signal sig_165:std_logic;
signal sig_166:std_logic;
signal sig_167:std_logic;
signal sig_168:std_logic;
signal sig_169:std_logic;
signal sig_170:std_logic;
signal sig_171:std_logic;
signal sig_5:std_logic_vector(1 downto 0);
signal sig_7:std_logic_vector(1 downto 0);
signal sig_9:std_logic_vector(1 downto 0);
signal sig_39:std_logic_vector(1 downto 0);
signal sig_41:std_logic_vector(1 downto 0);
signal sig_45:std_logic_vector(1 downto 0);
signal sig_46:std_logic_vector(1 downto 0);
signal sig_47:std_logic_vector(1 downto 0);
signal sig_48:std_logic_vector(1 downto 0);
signal sig_49:std_logic_vector(1 downto 0);
signal sig_50:std_logic_vector(1 downto 0);
signal sig_51:std_logic_vector(1 downto 0);
signal sig_52:std_logic_vector(1 downto 0);
signal sig_53:std_logic_vector(1 downto 0);
signal sig_54:std_logic_vector(1 downto 0);
signal sig_55:std_logic_vector(1 downto 0);
signal sig_63:std_logic_vector(1 downto 0);
signal sig_76:std_logic_vector(1 downto 0);
signal sig_77:std_logic_vector(1 downto 0);
signal CLK_Xv:std_logic;
signal CLK_Yv:std_logic;
signal CLK_Xp:std_logic;
signal CLK_Yp:std_logic;
signal CLK_Xfa:std_logic;
signal CLK_Yfa:std_logic;
signal CLK_Ga:std_logic;
signal CLK_Gb:std_logic;
signal CLK_Fa:std_logic;
signal CLK_Fb:std_logic;
signal CLK_Fc:std_logic;
signal CLK_Fd:std_logic;
signal CLK_TmpA:std_logic;
signal CLK_TmpB:std_logic;
signal CLK_ToMALU:std_logic;

--component map declaration
component wrapper_gf2m
   port(
      A:in std_logic_vector(162 downto 0);
      B:in std_logic_vector(162 downto 0);
      start:in std_logic;
      mode:in std_logic;
      plus_one:in std_logic;
      T:out std_logic_vector(162 downto 0);
      ready:out std_logic;
      RST : in std_logic;
      CLK : in std_logic
   );
end component;
type STATE_TYPE is (init1,init2,init3,init4,start,distort1,distort2,distort3,distort4,distort5,distort6,distort7,distort8,miller_init1,miller_init2,startloop1,ready1,ready2,dlambda1,dlambda2,dlambda3,dlambda4,s,alambda1,alambda2,alambda3,alambda4,alambda5,alambda6,alambda7,alambda8,alambda9,alambda10,alambda11,alambda12,alambda13,alambda14,alambda15,alambda16,alambda17,inv1,inv2,inv3,inv4,inv5,inv6,inv7,inv8,inv9,inv10,inv11,inv12,inv13,inv14,inv15,inv16,inv17,inv18,inv19,inv20,inv21,inv22,inv23,inv24,inv25,inv26,inv27,inv28,inv29,inv30,inv31,inv32,inv33,inv34,inv35,inv36,inv37,inv38,inv39,inv40,inv41,inv42,inv43,inv44,inv45,inv46,inv47,inv48,inv49,inv50,inv51,inv52,inv53,inv54,coord1,coord2,coord3,coord4,coord5,coord6,coord7,coord8,coord9,coord10,coord11,coord12,coord13,coord14,coord15,coord16,coord17,coord18,coord19,coord20,coord21,coord22,coord23,coord24,coord25,coord26,coord27,coord28,coord29,coord30,coord31,coord32,coord33,coord34,coord35,updatef1,fsqrt1,fsqrt2,fsqrt3,fsqrt4,fsqrt5,fsqrt6,fsqrt7,fsqrt8,fsqrt9,fsqrt10,fsqrt11,fsqrt12,fsqrt13,fsqrt14,fsqrt15,fsqrt16,fsqrt17,fsqrt18,fsqrt19,fsqrt20,fsqrt21,fsqrt22,fsqrt23,fsqrt24,fsqrt25,fsqrt26,fsqrt27,fsqrt28,fsqrt29,fsqrt30,fsqrt31,fsqrt32,fg1,fg2,fg3,fg4,fg5,fg6,fg7,fg8,fg9,fg10,fg11,fg12,fg13,fg14,fg15,fg16,fg17,fg18,fg19,fg20,fg21,fg22,fg23,fg24,fg25,fg26,fg27,fg28,fg29,fg30,fg31,fg32,fg33,fg34,fg35,fg36,fg37,fg38,fg39,fg40,fg41,fg42,fg43,fg44,fg45,fg46,fg47,fg48,fg49,fg50,fg51,fg52,fg53,fg54,fg55,fg56,fg57,fg58,fg59,fg60,fg61,fg62,fg63,fg64,fg65,fg66,fg67,finalexp1,finalexp2,finalexp3,finalexp4,finalexp5,finalexp6,finalexp7,finalexp8,finalexp9,finalexp10,finalexp11,finalexp12,finalexp13,finalexp14,finalexp15,finalexp16,finalexp17,finalexp18,finalexp19,finalexp20,finalexp21,finalexp22,finalexp23,finalexp24,finalexp25,finalexp26,finalexp27,finalexp28,finalexp29,finalexp30,finalexp31,finalexp32,finalexp33,finalexp34,finalexp35,finalexp36,finalexp37,finalexp38,finalexp39,finalexp40,finalexp41,finalexp42,finalexp43,finalexp44,finalexp45,finalexp46,finalexp47,finalexp48,finalexp49,finalexp50,finalexp51,finalexp52,finalexp53,finalexp54,finalexp55,finalexp56,finalexp57,finalexp58,finalexp59,finalexp60,finalexp61,finalexp62,finalexp63,finalexp64,finalexp65,finalexp66,finalexp67,finalexp68,finalexp69,finalexp70,finalexp71,finalexp72,finalexp73,finalexp74,finalexp75,finalexp76,finalexp77,finalexp78,finalexp79,finalexp80,f4mpow1,f4mpow2,f4mpow3,f4mpow4,f4mpow5,f4mpow6,f4mpow7,f4mpow8,f4mpow9,f4mpow10,f4mpow11,f4mpow12,f4mpow13,f4mpow14,f4mpow15,f4mpow16,f4mpow17,f4mpow18,f4mpow19,f4mpow20,f4mpow21,f4mpow22,f4mpow23,f4mpow24,f4mpow25,f4mpow26,f4mpow27,f4mpow28,f4mpow29,f4mpow30,f4mpow31,f4mpow32,f4mpow33,f4mpow34,f4mpow35,f4mpow36,f4mpow37,f4mpow38,f4mpow39,f4mpow40,f4mpow41,f4mpow42,f4mpow43,f4mpow44,f4mpow45,f4mpow46,f4mpow47,f4mpow48,f4mpow49,f4mpow50,f4mpow51,f4mpow52,f4mpow53,f4mpow54,f4mpow55,f4mpow56,f4mpow57,f4mpow58,f4mpow59,f4mpow60,f4mpow61,f4mpow62,f4mpow47fix,f4msqrt1,f4msqrt2,f4msqrt3,f4msqrt4,f4msqrt5,f4msqrt6,f4msqrt7,f4msqrt8,f4msqrt9,f4msqrt10,f4msqrt11,f4msqrt12,f4msqrt13,f4msqrt14,f4msqrt15,f4msqrt16,f4msqrt17,f4msqrt18,f4msqrt19,f4msqrt20,f4msqrt21,f4msqrt22,f4msqrt23,f4msqrt24,f4msqrt25,f4msqrt26,f4msqrt27,f4msqrt28,f4msqrt29,f4msqrt30,f4msqrt31,f4msqrt32,f4msqrt27fix,f4mmult1,f4mmult2,f4mmult3,f4mmult4,f4mmult5,f4mmult6,f4mmult7,f4mmult8,f4mmult9,f4mmult10,f4mmult11,f4mmult12,f4mmult13,f4mmult14,f4mmult15,f4mmult16,f4mmult17,f4mmult18,f4mmult19,f4mmult20,f4mmult21,f4mmult22,f4mmult23,f4mmult24,f4mmult25,f4mmult26,f4mmult27,f4mmult28,f4mmult29,f4mmult30,f4mmult31,f4mmult32,f4mmult33,f4mmult34,f4mmult35,f4mmult36,f4mmult37,f4mmult38,f4mmult39,f4mmult40,f4mmult41,f4mmult42,f4mmult43,f4mmult44,f4mmult45,f4mmult46,f4mmult47,f4mmult48,f4mmult49,f4mmult50,f4mmult51,f4mmult52,f4mmult53,f4mmult54,f4mmult55,f4mmult56,f4mmult57,f4mmult58,f4mmult59,f4mmult60,f4mmult61,f4mmult62,f4mmult63,f4mmult64,f4mmult65,f4mmult66,f4mmult67,f4mmult68,f4mmult69,f4mmult70,f4mmult71,f4mmult72,f4mmult73,f4mmult74,f4mmult75,f4mmult76,f4mmult77,f4mmult78,f4mmult79,f4mmult80,f4mmult81,f4mmult82,f4mmult83,f4mmult84,f4mmult85,f4mmult86,f4mmult87,f4mmult88,f4mmult89,f4mmult90,f4mmult91,f4mmult92,f4mmult93,f4mmult94,f4mmult95,f4mmult96,f4mmfix1,f4mmfix2,f4mmfix3,f4mmfix4,f4mmfix5,f2mmult1,f2mmult2,f2mmult3,f2mmult4,f2mmult5,f2mmult6,f2mmult7,f2mmult8,f2mmult9,f2mmult10,f2mmult11,f2mmult12,f2mmult13,f2mmult14,f2mmult15,f2mmult16,f2mmult17,f2mmult18,f2mmult19,f2mmult20,f2mmult21,f2mmult22,f2mmult23,f2mmult24,f2mmult25,f2mmult26,f2mmult27,f2mmult28,f2mmult29,f2minv1,f2minv2,f2minv3,f2minv4,f2minv5,f2minv6,f2minv7,f2minv8,f2minv9,f2minv10,f2minv11,f2minv12,f2minv13,f2minv14,f2minv15,f2minv16,f2minv17,f2minv18,f2minv19);
signal STATE:STATE_TYPE;
type CONTROL is (do_alwaysset_not_readyMALU_idleidle_ToMALUupdate_Xv_from_Inputidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_regs
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Inputidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Inputupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Inputupdate_Yv_from_Xvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_Inputupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysset_readyreset_counter_miscMALU_idleidle_regs
, do_alwaysready_regsMALU_idle
, do_alwaysMALU_addidle_regs
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleunset_addreset_Freset_counter_milleridle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_regsdec_counter_miller
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_mult_plus_oneidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaupdate_Gb_from_Faupdate_Fa_from_Fbupdate_Fb_from_Fcupdate_Fc_from_Fdidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_regsset_add
, do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaupdate_Gb_from_Faupdate_Fa_from_Fbupdate_Fb_from_Fcupdate_Fc_from_Fdidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_Fdupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysreset_counter_miscMALU_idleupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_multidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleidle_regsreset_counter_misc
, do_alwaysinc_counter_miscMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_add_plus_oneidle_ToMALUupdate_Xv_from_TmpBidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Gbupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xvupdate_Xp_from_Yvidle_Ypupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaupdate_Gb_from_Gaidle_Faidle_Fbupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_multupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_multupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Fcupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv
, do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_multidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_Fdupdate_TmpB_from_TmpA
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaupdate_Ga_from_Gbupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_Xv
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_TmpBidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaupdate_Yfa_from_Gaupdate_Ga_from_Gbidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_TmpAidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaupdate_Yfa_from_Gaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB
, unset_adddo_alwaysMALU_idleidle_regs
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_multupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Fcupdate_Fc_from_Fdupdate_Fd_from_TmpAidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBidle_TmpB
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Ypidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpupdate_Yp_from_Xpupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Ypupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaupdate_Yfa_from_Xfaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaupdate_Ga_from_Yfaupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaupdate_Ga_from_Gbupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaupdate_Gb_from_Gaupdate_Fa_from_Gbupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Gbupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaupdate_Gb_from_Faupdate_Fa_from_Gbidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaupdate_Ga_from_Gbupdate_Gb_from_Gaupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaupdate_Yfa_from_Gaupdate_Ga_from_Yfaupdate_Gb_from_Faupdate_Fa_from_Gbidle_Fbupdate_Fc_from_Fbidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaupdate_Ga_from_Gbupdate_Gb_from_Gaupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcupdate_Fd_from_Fcidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faupdate_Fc_from_Fbidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xfaidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Ypidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaupdate_Ga_from_Gbupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaupdate_Ga_from_Gbupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xfaidle_Xfaupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xfaidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA
, do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaupdate_Yfa_from_Xfaupdate_Ga_from_Yfaupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaupdate_Ga_from_Gbupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA
, do_alwaysinc_counter_miscMALU_idleidle_regs
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_Fdupdate_TmpB_from_TmpA
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Ypidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_Xv
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_Xv
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Yfaupdate_Yfa_from_Gaupdate_Ga_from_Gbidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_TmpBupdate_Yv_from_Xvupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaupdate_Yfa_from_Gaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Ypupdate_Yp_from_Xpupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_TmpBidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Fcupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaupdate_Gb_from_Faupdate_Fa_from_Fbupdate_Fb_from_Faupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAupdate_TmpB_from_TmpA
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbidle_Fdupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_Fcidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Faupdate_Fc_from_Fbidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB
, do_alwaysMALU_multidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcidle_TmpAidle_TmpB
, do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_addidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA
, do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Ypidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA
, do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
, do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaupdate_Gb_from_Gaupdate_Fa_from_Gbupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaupdate_Gb_from_Gaupdate_Fa_from_Gbupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA
, do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_multupdate_ToMALU_from_Xvupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB
, do_alwaysMALU_multupdate_ToMALU_from_Xvupdate_Xv_from_Yvupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv
);
signal cmd : CONTROL;


begin


   --portmap
   label_wrapper_gf2m : wrapper_gf2m port map (
         A => sig_MALU_A,
         B => sig_MALU_B,
         start => sig_MALU_start,
         mode => sig_MALU_mode,
         plus_one => sig_MALU_plus_one,
         T => sig_MALU_result,
         ready => sig_MALU_ready,
         RST => RST,
         CLK => CLK
      );
   --register updates
   dpREG: process (CLK,RST,CLK_Xv,CLK_Yv,CLK_Xp,CLK_Yp,CLK_Xfa,CLK_Yfa,CLK_Ga,CLK_Gb,CLK_Fa,CLK_Fb,CLK_Fc,CLK_Fd,CLK_TmpA,CLK_TmpB,CLK_ToMALU)
      begin
         if (RST = '1') then
            reg_counter_miller <= (others=>'0');
            reg_counter_misc <= (others=>'0');
            reg_add <= '0';
            reg_start <= '0';
            reg_next <= '0';
            reg_ready <= '0';
         elsif CLK' event and CLK = '1' then
            reg_MALU_ready <= reg_MALU_ready_wire;
            reg_counter_miller <= reg_counter_miller_wire;
            reg_counter_misc <= reg_counter_misc_wire;
            reg_add <= reg_add_wire;
            reg_start <= reg_start_wire;
            reg_next <= reg_next_wire;
            reg_ready <= reg_ready_wire;
	 end if;
   end process dpREG;

   process (CLK_Xv)
      begin
	 if CLK_Xv' event and CLK_Xv = '1' then
            reg_Xv <= reg_Xv_wire;
	 end if;	 
   end process;

   process (CLK_Yv)
      begin
	 if CLK_Yv' event and CLK_Yv = '1' then
            reg_Yv <= reg_Yv_wire;
	 end if;
   end process;

   process (CLK_Xp)
      begin
	 if CLK_Xp' event and CLK_Xp = '1' then
            reg_Xp <= reg_Xp_wire;
	 end if;
   end process;

   process (CLK_Yp)
      begin
	 if CLK_Yp' event and CLK_Yp = '1' then
            reg_Yp <= reg_Yp_wire;
	 end if;
   end process;

   process (CLK_Xfa)
      begin
	 if CLK_Xfa' event and CLK_Xfa = '1' then
            reg_Xfa <= reg_Xfa_wire;
	 end if;
   end process;

   process (CLK_Yfa)
      begin
	 if CLK_Yfa' event and CLK_Yfa = '1' then
            reg_Yfa <= reg_Yfa_wire;
	 end if;
   end process;

   process (CLK_Ga)
      begin
	 if CLK_Ga' event and CLK_Ga = '1' then
            reg_Ga <= reg_Ga_wire;
	 end if;
   end process;

   process (CLK_Gb)
      begin
	 if CLK_Gb' event and CLK_Gb = '1' then
            reg_Gb <= reg_Gb_wire;
	 end if;
   end process;

   process (CLK_Fa)
      begin
	 if CLK_Fa' event and CLK_Fa = '1' then
            reg_Fa <= reg_Fa_wire;
	 end if;
   end process;

   process (CLK_Fb)
      begin
	 if CLK_Fb' event and CLK_Fb = '1' then
            reg_Fb <= reg_Fb_wire;
	 end if;
   end process;

   process (CLK_Fc)
      begin
	 if CLK_Fc' event and CLK_Fc = '1' then
            reg_Fc <= reg_Fc_wire;
	 end if;
   end process;

   process (CLK_Fd)
      begin
	 if CLK_Fd' event and CLK_Fd = '1' then
            reg_Fd <= reg_Fd_wire;
	 end if;
   end process;

   process (CLK_TmpA)
      begin
	 if CLK_TmpA' event and CLK_TmpA = '1' then
            reg_TmpA <= reg_TmpA_wire;
	 end if;
   end process;

   process (CLK_TmpB)
      begin
	 if CLK_TmpB' event and CLK_TmpB = '1' then
            reg_TmpB <= reg_TmpB_wire;
	 end if;
   end process;

   process (CLK_ToMALU)
      begin
	 if CLK_ToMALU' event and CLK_ToMALU = '1' then
            reg_ToMALU <= reg_ToMALU_wire;
         end if;
      end process;


   --combinational logics
   dpCMB: process (reg_Xv,reg_Yv,reg_Xp,reg_Yp,reg_Xfa,reg_Yfa,reg_Ga,reg_Gb,reg_Fa,reg_Fb
,reg_Fc,reg_Fd,reg_TmpA,reg_TmpB,reg_ToMALU,reg_MALU_ready,reg_counter_miller,reg_counter_misc,reg_add,reg_start
,reg_next,reg_ready,sig_MALU_A,sig_MALU_B,sig_MALU_start,sig_MALU_mode,sig_MALU_plus_one,sig_MALU_result,sig_MALU_ready,sig_en_Xv
,sig_en_Yv,sig_en_Xp,sig_en_Yp,sig_en_Xfa,sig_en_Yfa,sig_en_Ga,sig_en_Gb,sig_en_Fa,sig_en_Fb,sig_en_Fc
,sig_en_Fd,sig_en_TmpA,sig_en_TmpB,sig_en_ToMALU,sig_sel_Xv,sig_sel_Yv,sig_sel_Xp,sig_sel_Yp,sig_sel_Xfa,sig_sel_Yfa
,sig_sel_Ga,sig_sel_Gb,sig_sel_Fa,sig_sel_Fb,sig_sel_Fc,sig_sel_Fd,sig_sel_TmpA,sig_sel_TmpB,sig_sel_ToMALU,sig_to_Xv
,sig_to_Yv,sig_to_Xp,sig_to_Yp,sig_to_Xfa,sig_to_Yfa,sig_to_Ga,sig_to_Gb,sig_to_Fa,sig_to_Fb,sig_to_Fc
,sig_to_Fd,sig_to_TmpA,sig_to_TmpB,sig_to_ToMALU,sig_from_Xv,sig_from_Yv,sig_from_Xp,sig_from_Yp,sig_from_Xfa,sig_from_Yfa
,sig_from_Ga,sig_from_Gb,sig_from_Fa,sig_from_Fb,sig_from_Fc,sig_from_Fd,sig_from_TmpA,sig_from_TmpB,sig_from_ToMALU,sig_from_ToMALUShift
,sig_from_Input,sig_0,sig_1,sig_2,sig_3,sig_4,sig_6,sig_8,sig_10,sig_11
,sig_12,sig_13,sig_14,sig_15,sig_16,sig_17,sig_18,sig_19,sig_20,sig_21
,sig_22,sig_23,sig_24,sig_25,sig_26,sig_27,sig_28,sig_29,sig_30,sig_31
,sig_32,sig_33,sig_34,sig_35,sig_36,sig_37,sig_38,sig_40,sig_42,sig_43
,sig_44,sig_56,sig_57,sig_58,sig_59,sig_60,sig_61,sig_62,sig_64,sig_65
,sig_66,sig_67,sig_68,sig_69,sig_70,sig_71,sig_72,sig_73,sig_74,sig_75
,ready_int,output_int,sig_en_out_Xv_int,sig_en_out_Yv_int,sig_en_out_Xp_int,sig_en_out_Yp_int,sig_en_out_Xfa_int,sig_en_out_Yfa_int,sig_en_out_Ga_int,sig_en_out_Gb_int
,sig_en_out_Fa_int,sig_en_out_Fb_int,sig_en_out_Fc_int,sig_en_out_Fd_int,sig_en_out_TmpA_int,sig_en_out_TmpB_int,sig_en_out_ToMALU_int,input,start_in,next_in
,cmd,STATE)
      begin
         reg_Xv_wire <= reg_Xv;
         reg_Yv_wire <= reg_Yv;
         reg_Xp_wire <= reg_Xp;
         reg_Yp_wire <= reg_Yp;
         reg_Xfa_wire <= reg_Xfa;
         reg_Yfa_wire <= reg_Yfa;
         reg_Ga_wire <= reg_Ga;
         reg_Gb_wire <= reg_Gb;
         reg_Fa_wire <= reg_Fa;
         reg_Fb_wire <= reg_Fb;
         reg_Fc_wire <= reg_Fc;
         reg_Fd_wire <= reg_Fd;
         reg_TmpA_wire <= reg_TmpA;
         reg_TmpB_wire <= reg_TmpB;
         reg_ToMALU_wire <= reg_ToMALU;
         reg_MALU_ready_wire <= reg_MALU_ready;
         reg_counter_miller_wire <= reg_counter_miller;
         reg_counter_misc_wire <= reg_counter_misc;
         reg_add_wire <= reg_add;
         reg_start_wire <= reg_start;
         reg_next_wire <= reg_next;
         reg_ready_wire <= reg_ready;
         sig_MALU_A <= (others=>'0');
         sig_MALU_B <= (others=>'0');
         sig_MALU_start <= '0';
         sig_MALU_mode <= '0';
         sig_MALU_plus_one <= '0';
         sig_en_Xv <= '0';
         sig_en_Yv <= '0';
         sig_en_Xp <= '0';
         sig_en_Yp <= '0';
         sig_en_Xfa <= '0';
         sig_en_Yfa <= '0';
         sig_en_Ga <= '0';
         sig_en_Gb <= '0';
         sig_en_Fa <= '0';
         sig_en_Fb <= '0';
         sig_en_Fc <= '0';
         sig_en_Fd <= '0';
         sig_en_TmpA <= '0';
         sig_en_TmpB <= '0';
         sig_en_ToMALU <= '0';
         sig_sel_Xv <= (others=>'0');
         sig_sel_Yv <= '0';
         sig_sel_Xp <= '0';
         sig_sel_Yp <= '0';
         sig_sel_Xfa <= '0';
         sig_sel_Yfa <= '0';
         sig_sel_Ga <= '0';
         sig_sel_Gb <= '0';
         sig_sel_Fa <= '0';
         sig_sel_Fb <= '0';
         sig_sel_Fc <= '0';
         sig_sel_Fd <= '0';
         sig_sel_TmpA <= '0';
         sig_sel_TmpB <= '0';
         sig_sel_ToMALU <= (others=>'0');
         sig_to_Xv <= (others=>'0');
         sig_to_Yv <= (others=>'0');
         sig_to_Xp <= (others=>'0');
         sig_to_Yp <= (others=>'0');
         sig_to_Xfa <= (others=>'0');
         sig_to_Yfa <= (others=>'0');
         sig_to_Ga <= (others=>'0');
         sig_to_Gb <= (others=>'0');
         sig_to_Fa <= (others=>'0');
         sig_to_Fb <= (others=>'0');
         sig_to_Fc <= (others=>'0');
         sig_to_Fd <= (others=>'0');
         sig_to_TmpA <= (others=>'0');
         sig_to_TmpB <= (others=>'0');
         sig_to_ToMALU <= (others=>'0');
         sig_from_Xv <= (others=>'0');
         sig_from_Yv <= (others=>'0');
         sig_from_Xp <= (others=>'0');
         sig_from_Yp <= (others=>'0');
         sig_from_Xfa <= (others=>'0');
         sig_from_Yfa <= (others=>'0');
         sig_from_Ga <= (others=>'0');
         sig_from_Gb <= (others=>'0');
         sig_from_Fa <= (others=>'0');
         sig_from_Fb <= (others=>'0');
         sig_from_Fc <= (others=>'0');
         sig_from_Fd <= (others=>'0');
         sig_from_TmpA <= (others=>'0');
         sig_from_TmpB <= (others=>'0');
         sig_from_ToMALU <= (others=>'0');
         sig_from_ToMALUShift <= (others=>'0');
         sig_from_Input <= (others=>'0');
         sig_0 <= '0';
         sig_1 <= (others=>'0');
         sig_2 <= (others=>'0');
         sig_3 <= '0';
         sig_4 <= (others=>'0');
         sig_6 <= '0';
         sig_8 <= '0';
         sig_10 <= '0';
         sig_11 <= (others=>'0');
         sig_12 <= (others=>'0');
         sig_13 <= '0';
         sig_14 <= (others=>'0');
         sig_15 <= '0';
         sig_16 <= (others=>'0');
         sig_17 <= '0';
         sig_18 <= (others=>'0');
         sig_19 <= '0';
         sig_20 <= (others=>'0');
         sig_21 <= '0';
         sig_22 <= (others=>'0');
         sig_23 <= '0';
         sig_24 <= (others=>'0');
         sig_25 <= '0';
         sig_26 <= (others=>'0');
         sig_27 <= '0';
         sig_28 <= (others=>'0');
         sig_29 <= '0';
         sig_30 <= (others=>'0');
         sig_31 <= '0';
         sig_32 <= (others=>'0');
         sig_33 <= '0';
         sig_34 <= (others=>'0');
         sig_35 <= '0';
         sig_36 <= (others=>'0');
         sig_37 <= '0';
         sig_38 <= (others=>'0');
         sig_40 <= '0';
         sig_42 <= '0';
         sig_43 <= (others=>'0');
         sig_44 <= (others=>'0');
         sig_56 <= (others=>'0');
         sig_57 <= (others=>'0');
         sig_58 <= '0';
         sig_59 <= '0';
         sig_60 <= '0';
         sig_61 <= (others=>'0');
         sig_62 <= (others=>'0');
         sig_64 <= '0';
         sig_65 <= '0';
         sig_66 <= '0';
         sig_67 <= (others=>'0');
         sig_68 <= '0';
         sig_69 <= '0';
         sig_70 <= '0';
         sig_71 <= (others=>'0');
         sig_72 <= '0';
         sig_73 <= '0';
         sig_74 <= '0';
         sig_75 <= (others=>'0');
         ready_int <= '0';
         output_int <= (others=>'0');
         sig_en_out_Xv_int <= '0';
         sig_en_out_Yv_int <= '0';
         sig_en_out_Xp_int <= '0';
         sig_en_out_Yp_int <= '0';
         sig_en_out_Xfa_int <= '0';
         sig_en_out_Yfa_int <= '0';
         sig_en_out_Ga_int <= '0';
         sig_en_out_Gb_int <= '0';
         sig_en_out_Fa_int <= '0';
         sig_en_out_Fb_int <= '0';
         sig_en_out_Fc_int <= '0';
         sig_en_out_Fd_int <= '0';
         sig_en_out_TmpA_int <= '0';
         sig_en_out_TmpB_int <= '0';
         sig_en_out_ToMALU_int <= '0';
         sig_5 <= "10";
         sig_7 <= "11";
         sig_9 <= "00";
         sig_39 <= "00";
         sig_41 <= "01";
         sig_45 <= "00";
         sig_46 <= "00";
         sig_47 <= "00";
         sig_48 <= "00";
         sig_49 <= "00";
         sig_50 <= "01";
         sig_51 <= "11";
         sig_52 <= "11";
         sig_53 <= "10";
         sig_54 <= "01";
         sig_55 <= "00";
         sig_63 <= "01";
         sig_76 <= "00";
         sig_77 <= "00";
         output <= (others=>'0');
         ready <= '0';
         sig_en_out_Xv <= '0';
         sig_en_out_Yv <= '0';
         sig_en_out_Xp <= '0';
         sig_en_out_Yp <= '0';
         sig_en_out_Xfa <= '0';
         sig_en_out_Yfa <= '0';
         sig_en_out_Ga <= '0';
         sig_en_out_Gb <= '0';
         sig_en_out_Fa <= '0';
         sig_en_out_Fb <= '0';
         sig_en_out_Fc <= '0';
         sig_en_out_Fd <= '0';
         sig_en_out_TmpA <= '0';
         sig_en_out_TmpB <= '0';
         sig_en_out_ToMALU <= '0';



         case cmd is
            when do_alwaysset_not_readyMALU_idleidle_ToMALUupdate_Xv_from_Inputidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               reg_ready_wire <= '0';
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_52;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_regs =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_Xv <= '0';
               sig_en_Yv <= '0';
               sig_en_Xp <= '0';
               sig_en_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_en_Gb <= '0';
               sig_en_Fa <= '0';
               sig_en_Fb <= '0';
               sig_en_Fc <= '0';
               sig_en_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_Xv <= sig_45;
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '0';
               sig_sel_Yfa <= '0';
               sig_sel_Ga <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '0';
               sig_sel_ToMALU <= sig_46;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Inputidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_52;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Inputupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_52;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Inputupdate_Yv_from_Xvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_52;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_Inputupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_52;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysset_readyreset_counter_miscMALU_idleidle_regs =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               reg_ready_wire <= '1';
               reg_TmpB_wire <= conv_std_logic_vector(0,163);
               reg_counter_misc_wire <= conv_std_logic_vector(0,7);
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_Xv <= '0';
               sig_en_Yv <= '0';
               sig_en_Xp <= '0';
               sig_en_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_en_Gb <= '0';
               sig_en_Fa <= '0';
               sig_en_Fb <= '0';
               sig_en_Fc <= '0';
               sig_en_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_Xv <= sig_45;
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '0';
               sig_sel_Yfa <= '0';
               sig_sel_Ga <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '0';
               sig_sel_ToMALU <= sig_46;
            when do_alwaysready_regsMALU_idle =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               if (next_in = '1') then
                  sig_58 <= '1';
               else
                  sig_58 <= '0';
               end if;
               if (reg_next = '0') then
                  sig_59 <= '1';
               else
                  sig_59 <= '0';
               end if;
               sig_60 <= sig_58 and sig_59;
               sig_61 <= unsigned(reg_counter_misc) + unsigned(conv_std_logic_vector(1,7));
               if (sig_60 = '1') then
                  sig_62 <= sig_61;
               else
                  sig_62 <= reg_counter_misc;
               end if;
               sig_en_Xv <= '1';
               sig_en_Yv <= '1';
               sig_en_Xp <= '1';
               sig_sel_Xv <= sig_63;
               sig_sel_Yv <= '1';
               sig_sel_Xp <= '1';
               if (next_in = '1') then
                  sig_64 <= '1';
               else
                  sig_64 <= '0';
               end if;
               if (reg_next = '0') then
                  sig_65 <= '1';
               else
                  sig_65 <= '0';
               end if;
               sig_66 <= sig_64 and sig_65;
               if (sig_66 = '1') then
                  sig_67 <= sig_to_Xv;
               else
                  sig_67 <= reg_Xv;
               end if;
               if (next_in = '1') then
                  sig_68 <= '1';
               else
                  sig_68 <= '0';
               end if;
               if (reg_next = '0') then
                  sig_69 <= '1';
               else
                  sig_69 <= '0';
               end if;
               sig_70 <= sig_68 and sig_69;
               if (sig_70 = '1') then
                  sig_71 <= sig_to_Yv;
               else
                  sig_71 <= reg_Yv;
               end if;
               if (next_in = '1') then
                  sig_72 <= '1';
               else
                  sig_72 <= '0';
               end if;
               if (reg_next = '0') then
                  sig_73 <= '1';
               else
                  sig_73 <= '0';
               end if;
               sig_74 <= sig_72 and sig_73;
               if (sig_74 = '1') then
                  sig_75 <= sig_to_Xp;
               else
                  sig_75 <= reg_Xp;
               end if;
               sig_en_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_en_Gb <= '0';
               sig_en_Fa <= '0';
               sig_en_Fb <= '0';
               sig_en_Fc <= '0';
               sig_en_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_en_ToMALU <= sig_76(0);
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '0';
               sig_sel_Yfa <= '0';
               sig_sel_Ga <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '0';
               sig_sel_ToMALU <= sig_77;
               reg_counter_misc_wire <= sig_62;
               reg_Xv_wire <= sig_67;
               reg_Yv_wire <= sig_71;
               reg_Xp_wire <= sig_75;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
            when do_alwaysMALU_addidle_regs =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_Xv <= '0';
               sig_en_Yv <= '0';
               sig_en_Xp <= '0';
               sig_en_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_en_Gb <= '0';
               sig_en_Fa <= '0';
               sig_en_Fb <= '0';
               sig_en_Fc <= '0';
               sig_en_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_Xv <= sig_45;
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '0';
               sig_sel_Yfa <= '0';
               sig_sel_Ga <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '0';
               sig_sel_ToMALU <= sig_46;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleunset_addreset_Freset_counter_milleridle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               reg_add_wire <= '0';
               reg_Fa_wire <= conv_std_logic_vector(1,163);
               reg_Fb_wire <= conv_std_logic_vector(0,163);
               reg_Fc_wire <= conv_std_logic_vector(0,163);
               reg_Fd_wire <= conv_std_logic_vector(0,163);
               reg_counter_miller_wire <= conv_std_logic_vector(163,8);
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_regsdec_counter_miller =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_Xv <= '0';
               sig_en_Yv <= '0';
               sig_en_Xp <= '0';
               sig_en_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_en_Gb <= '0';
               sig_en_Fa <= '0';
               sig_en_Fb <= '0';
               sig_en_Fc <= '0';
               sig_en_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_Xv <= sig_45;
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '0';
               sig_sel_Yfa <= '0';
               sig_sel_Ga <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '0';
               sig_sel_ToMALU <= sig_46;
               sig_56 <= unsigned(reg_counter_miller) - unsigned(conv_std_logic_vector(1,8));
               reg_counter_miller_wire <= sig_56;
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_mult_plus_oneidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '1';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_51;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaupdate_Gb_from_Faupdate_Fa_from_Fbupdate_Fb_from_Fcupdate_Fc_from_Fdidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '0';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_sel_Gb <= '1';
               sig_en_Gb <= '1';
               reg_Gb_wire <= sig_to_Gb;
               sig_sel_Fa <= '1';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_regsset_add =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_Xv <= '0';
               sig_en_Yv <= '0';
               sig_en_Xp <= '0';
               sig_en_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_en_Gb <= '0';
               sig_en_Fa <= '0';
               sig_en_Fb <= '0';
               sig_en_Fc <= '0';
               sig_en_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_Xv <= sig_45;
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '0';
               sig_sel_Yfa <= '0';
               sig_sel_Ga <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '0';
               sig_sel_ToMALU <= sig_46;
               reg_add_wire <= '1';
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaupdate_Gb_from_Faupdate_Fa_from_Fbupdate_Fb_from_Fcupdate_Fc_from_Fdidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_sel_Gb <= '1';
               sig_en_Gb <= '1';
               reg_Gb_wire <= sig_to_Gb;
               sig_sel_Fa <= '1';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_Fdupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '0';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysreset_counter_miscMALU_idleupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               reg_counter_misc_wire <= conv_std_logic_vector(0,7);
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_multidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_regsreset_counter_misc =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_Xv <= '0';
               sig_en_Yv <= '0';
               sig_en_Xp <= '0';
               sig_en_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_en_Gb <= '0';
               sig_en_Fa <= '0';
               sig_en_Fb <= '0';
               sig_en_Fc <= '0';
               sig_en_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_Xv <= sig_45;
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '0';
               sig_sel_Yfa <= '0';
               sig_sel_Ga <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '0';
               sig_sel_ToMALU <= sig_46;
               reg_counter_misc_wire <= conv_std_logic_vector(0,7);
            when do_alwaysinc_counter_miscMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_57 <= unsigned(reg_counter_misc) + unsigned(conv_std_logic_vector(1,7));
               reg_counter_misc_wire <= sig_57;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '1';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '0';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_add_plus_oneidle_ToMALUupdate_Xv_from_TmpBidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '1';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Gbupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xvupdate_Xp_from_Yvidle_Ypupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaupdate_Gb_from_Gaidle_Faidle_Fbupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '0';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_sel_Gb <= '0';
               sig_en_Gb <= '1';
               reg_Gb_wire <= sig_to_Gb;
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Fcupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '1';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '1';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '1';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '1';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_multidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_Fdupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '1';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '0';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '1';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaupdate_Ga_from_Gbupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '1';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_sel_Gb <= '0';
               sig_en_Gb <= '1';
               reg_Gb_wire <= sig_to_Gb;
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_TmpBidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_sel_Yfa <= '1';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '0';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaupdate_Yfa_from_Gaupdate_Ga_from_Gbidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_TmpAidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '1';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '1';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaupdate_Yfa_from_Gaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '1';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when unset_adddo_alwaysMALU_idleidle_regs =>
               reg_add_wire <= '0';
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_Xv <= '0';
               sig_en_Yv <= '0';
               sig_en_Xp <= '0';
               sig_en_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_en_Gb <= '0';
               sig_en_Fa <= '0';
               sig_en_Fb <= '0';
               sig_en_Fc <= '0';
               sig_en_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_Xv <= sig_45;
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '0';
               sig_sel_Yfa <= '0';
               sig_sel_Ga <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '0';
               sig_sel_ToMALU <= sig_46;
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Fcupdate_Fc_from_Fdupdate_Fd_from_TmpAidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '1';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Ypidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpupdate_Yp_from_Xpupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '1';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Ypupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaupdate_Yfa_from_Xfaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '0';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaupdate_Ga_from_Yfaupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_sel_Ga <= '0';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_sel_Gb <= '0';
               sig_en_Gb <= '1';
               reg_Gb_wire <= sig_to_Gb;
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaupdate_Ga_from_Gbupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_sel_Ga <= '1';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_sel_Gb <= '0';
               sig_en_Gb <= '1';
               reg_Gb_wire <= sig_to_Gb;
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaupdate_Gb_from_Gaupdate_Fa_from_Gbupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_sel_Gb <= '0';
               sig_en_Gb <= '1';
               reg_Gb_wire <= sig_to_Gb;
               sig_sel_Fa <= '0';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Gbupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaupdate_Gb_from_Faupdate_Fa_from_Gbidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_sel_Gb <= '1';
               sig_en_Gb <= '1';
               reg_Gb_wire <= sig_to_Gb;
               sig_sel_Fa <= '0';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaupdate_Ga_from_Gbupdate_Gb_from_Gaupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_sel_Ga <= '1';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_sel_Gb <= '0';
               sig_en_Gb <= '1';
               reg_Gb_wire <= sig_to_Gb;
               sig_sel_Fa <= '1';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaupdate_Yfa_from_Gaupdate_Ga_from_Yfaupdate_Gb_from_Faupdate_Fa_from_Gbidle_Fbupdate_Fc_from_Fbidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_sel_Yfa <= '1';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '0';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_sel_Gb <= '1';
               sig_en_Gb <= '1';
               reg_Gb_wire <= sig_to_Gb;
               sig_sel_Fa <= '0';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaupdate_Ga_from_Gbupdate_Gb_from_Gaupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcupdate_Fd_from_Fcidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '1';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_sel_Gb <= '0';
               sig_en_Gb <= '1';
               reg_Gb_wire <= sig_to_Gb;
               sig_sel_Fa <= '1';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faupdate_Fc_from_Fbidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_sel_Yfa <= '1';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '0';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '1';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xfaidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Ypidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaupdate_Ga_from_Gbupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_sel_Ga <= '1';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_sel_Gb <= '0';
               sig_en_Gb <= '1';
               reg_Gb_wire <= sig_to_Gb;
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_sel_Yfa <= '1';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '0';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaupdate_Ga_from_Gbupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '1';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_sel_Gb <= '0';
               sig_en_Gb <= '1';
               reg_Gb_wire <= sig_to_Gb;
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xfaidle_Xfaupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_sel_Yfa <= '1';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '0';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xfaidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '0';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '0';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaupdate_Yfa_from_Xfaupdate_Ga_from_Yfaupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '0';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_sel_Gb <= '0';
               sig_en_Gb <= '1';
               reg_Gb_wire <= sig_to_Gb;
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_sel_Yfa <= '1';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '0';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaupdate_Ga_from_Gbupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_sel_Ga <= '1';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_sel_Gb <= '0';
               sig_en_Gb <= '1';
               reg_Gb_wire <= sig_to_Gb;
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysinc_counter_miscMALU_idleidle_regs =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_57 <= unsigned(reg_counter_misc) + unsigned(conv_std_logic_vector(1,7));
               reg_counter_misc_wire <= sig_57;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_Xv <= '0';
               sig_en_Yv <= '0';
               sig_en_Xp <= '0';
               sig_en_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_en_Gb <= '0';
               sig_en_Fa <= '0';
               sig_en_Fb <= '0';
               sig_en_Fc <= '0';
               sig_en_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_Xv <= sig_45;
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '0';
               sig_sel_Yfa <= '0';
               sig_sel_Ga <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '0';
               sig_sel_ToMALU <= sig_46;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_Fdupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Ypidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Yfaupdate_Yfa_from_Gaupdate_Ga_from_Gbidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '1';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '1';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_TmpBupdate_Yv_from_Xvupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaupdate_Yfa_from_Gaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '1';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Ypupdate_Yp_from_Xpupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_TmpBidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Fcupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '1';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaupdate_Gb_from_Faupdate_Fa_from_Fbupdate_Fb_from_Faupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_sel_Gb <= '1';
               sig_en_Gb <= '1';
               reg_Gb_wire <= sig_to_Gb;
               sig_sel_Fa <= '1';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '1';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbidle_Fdupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_Fcidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Faupdate_Fc_from_Fbidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_sel_Fc <= '1';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_sel_Fa <= '1';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '1';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '1';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '1';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_addidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '1';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Ypidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_50;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_sel_TmpA <= '1';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '1';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaupdate_Gb_from_Gaupdate_Fa_from_Gbupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_sel_Yv <= '0';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '0';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_sel_Gb <= '0';
               sig_en_Gb <= '1';
               reg_Gb_wire <= sig_to_Gb;
               sig_sel_Fa <= '0';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaupdate_Gb_from_Gaupdate_Fa_from_Gbupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_en_Xv <= '0';
               sig_sel_Xv <= sig_47;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_sel_Yp <= '0';
               sig_en_Yp <= '1';
               reg_Yp_wire <= sig_to_Yp;
               sig_sel_Xfa <= '0';
               sig_en_Xfa <= '1';
               reg_Xfa_wire <= sig_to_Xfa;
               sig_sel_Yfa <= '0';
               sig_en_Yfa <= '1';
               reg_Yfa_wire <= sig_to_Yfa;
               sig_sel_Ga <= '0';
               sig_en_Ga <= '1';
               reg_Ga_wire <= sig_to_Ga;
               sig_sel_Gb <= '0';
               sig_en_Gb <= '1';
               reg_Gb_wire <= sig_to_Gb;
               sig_sel_Fa <= '0';
               sig_en_Fa <= '1';
               reg_Fa_wire <= sig_to_Fa;
               sig_sel_Fb <= '0';
               sig_en_Fb <= '1';
               reg_Fb_wire <= sig_to_Fb;
               sig_sel_Fc <= '0';
               sig_en_Fc <= '1';
               reg_Fc_wire <= sig_to_Fc;
               sig_sel_Fd <= '0';
               sig_en_Fd <= '1';
               reg_Fd_wire <= sig_to_Fd;
               sig_sel_TmpA <= '0';
               sig_en_TmpA <= '1';
               reg_TmpA_wire <= sig_to_TmpA;
               sig_sel_TmpB <= '0';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '0';
               sig_MALU_mode <= '0';
               sig_MALU_plus_one <= '0';
               sig_en_ToMALU <= '0';
               sig_sel_ToMALU <= sig_48;
               sig_sel_Xv <= sig_53;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_sel_Xp <= '0';
               sig_en_Xp <= '1';
               reg_Xp_wire <= sig_to_Xp;
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multupdate_ToMALU_from_Xvupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_55;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_en_Yv <= '0';
               sig_sel_Yv <= '0';
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_en_TmpB <= '0';
               sig_sel_TmpB <= '0';
            when do_alwaysMALU_multupdate_ToMALU_from_Xvupdate_Xv_from_Yvupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv =>
               ready <= ready_int;
               if (reg_ready = '0') then
                  sig_0 <= '1';
               else
                  sig_0 <= '0';
               end if;
               if (sig_0 = '1') then
                  sig_1 <= conv_std_logic_vector(0,163);
               else
                  sig_1 <= sig_from_Xv;
               end if;
               output <= output_int;
               sig_MALU_A <= reg_ToMALU;
               sig_MALU_B <= reg_Xv;
               sig_en_out_Xv <= sig_en_out_Xv_int;
               sig_en_out_Yv <= sig_en_out_Yv_int;
               sig_en_out_Xp <= sig_en_out_Xp_int;
               sig_en_out_Yp <= sig_en_out_Yp_int;
               sig_en_out_Xfa <= sig_en_out_Xfa_int;
               sig_en_out_Yfa <= sig_en_out_Yfa_int;
               sig_en_out_Ga <= sig_en_out_Ga_int;
               sig_en_out_Gb <= sig_en_out_Gb_int;
               sig_en_out_Fa <= sig_en_out_Fa_int;
               sig_en_out_Fb <= sig_en_out_Fb_int;
               sig_en_out_Fc <= sig_en_out_Fc_int;
               sig_en_out_Fd <= sig_en_out_Fd_int;
               sig_en_out_TmpA <= sig_en_out_TmpA_int;
               sig_en_out_TmpB <= sig_en_out_TmpB_int;
               sig_en_out_ToMALU <= sig_en_out_ToMALU_int;
               sig_from_Xv <= reg_Xv;
               sig_from_Yv <= reg_Yv;
               sig_from_Xp <= reg_Xp;
               sig_from_Yp <= reg_Yp;
               sig_from_Xfa <= reg_Xfa;
               sig_from_Yfa <= reg_Yfa;
               sig_from_Ga <= reg_Ga;
               sig_from_Gb <= reg_Gb;
               sig_from_Fa <= reg_Fa;
               sig_from_Fb <= reg_Fb;
               sig_from_Fc <= reg_Fc;
               sig_from_Fd <= reg_Fd;
               sig_from_TmpA <= reg_TmpA;
               sig_from_TmpB <= reg_TmpB;
               sig_from_ToMALU <= reg_ToMALU;
               sig_2 <= conv_std_logic_vector(signed(reg_ToMALU(161 downto 0)),162);
               sig_3 <= reg_ToMALU(162);
               sig_4 <= sig_2 & sig_3;
               sig_from_ToMALUShift <= sig_4;
               sig_from_Input <= input;
               if (unsigned(sig_sel_Xv) = unsigned(sig_5)) then
                  sig_6 <= '1';
               else
                  sig_6 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_7)) then
                  sig_8 <= '1';
               else
                  sig_8 <= '0';
               end if;
               if (unsigned(sig_sel_Xv) = unsigned(sig_9)) then
                  sig_10 <= '1';
               else
                  sig_10 <= '0';
               end if;
               if (sig_10 = '1') then
                  sig_11 <= sig_from_TmpB;
               else
                  sig_11 <= sig_from_Yv;
               end if;
               if (sig_6 = '1') then
                  sig_12 <= sig_from_ToMALU;
               elsif (sig_8 = '1') then
                  sig_12 <= sig_from_Input;
               else
                  sig_12 <= sig_11;
               end if;
               sig_to_Xv <= sig_12;
               if (sig_sel_Yv = '0') then
                  sig_13 <= '1';
               else
                  sig_13 <= '0';
               end if;
               if (sig_13 = '1') then
                  sig_14 <= sig_from_Xv;
               else
                  sig_14 <= sig_from_Xp;
               end if;
               sig_to_Yv <= sig_14;
               if (sig_sel_Xp = '0') then
                  sig_15 <= '1';
               else
                  sig_15 <= '0';
               end if;
               if (sig_15 = '1') then
                  sig_16 <= sig_from_Yv;
               else
                  sig_16 <= sig_from_Yp;
               end if;
               sig_to_Xp <= sig_16;
               if (sig_sel_Yp = '0') then
                  sig_17 <= '1';
               else
                  sig_17 <= '0';
               end if;
               if (sig_17 = '1') then
                  sig_18 <= sig_from_Xp;
               else
                  sig_18 <= sig_from_Xfa;
               end if;
               sig_to_Yp <= sig_18;
               if (sig_sel_Xfa = '0') then
                  sig_19 <= '1';
               else
                  sig_19 <= '0';
               end if;
               if (sig_19 = '1') then
                  sig_20 <= sig_from_Yp;
               else
                  sig_20 <= sig_from_Yfa;
               end if;
               sig_to_Xfa <= sig_20;
               if (sig_sel_Yfa = '0') then
                  sig_21 <= '1';
               else
                  sig_21 <= '0';
               end if;
               if (sig_21 = '1') then
                  sig_22 <= sig_from_Xfa;
               else
                  sig_22 <= sig_from_Ga;
               end if;
               sig_to_Yfa <= sig_22;
               if (sig_sel_Ga = '0') then
                  sig_23 <= '1';
               else
                  sig_23 <= '0';
               end if;
               if (sig_23 = '1') then
                  sig_24 <= sig_from_Yfa;
               else
                  sig_24 <= sig_from_Gb;
               end if;
               sig_to_Ga <= sig_24;
               if (sig_sel_Gb = '0') then
                  sig_25 <= '1';
               else
                  sig_25 <= '0';
               end if;
               if (sig_25 = '1') then
                  sig_26 <= sig_from_Ga;
               else
                  sig_26 <= sig_from_Fa;
               end if;
               sig_to_Gb <= sig_26;
               if (sig_sel_Fa = '0') then
                  sig_27 <= '1';
               else
                  sig_27 <= '0';
               end if;
               if (sig_27 = '1') then
                  sig_28 <= sig_from_Gb;
               else
                  sig_28 <= sig_from_Fb;
               end if;
               sig_to_Fa <= sig_28;
               if (sig_sel_Fb = '0') then
                  sig_29 <= '1';
               else
                  sig_29 <= '0';
               end if;
               if (sig_29 = '1') then
                  sig_30 <= sig_from_Fa;
               else
                  sig_30 <= sig_from_Fc;
               end if;
               sig_to_Fb <= sig_30;
               if (sig_sel_Fc = '0') then
                  sig_31 <= '1';
               else
                  sig_31 <= '0';
               end if;
               if (sig_31 = '1') then
                  sig_32 <= sig_from_Fb;
               else
                  sig_32 <= sig_from_Fd;
               end if;
               sig_to_Fc <= sig_32;
               if (sig_sel_Fd = '0') then
                  sig_33 <= '1';
               else
                  sig_33 <= '0';
               end if;
               if (sig_33 = '1') then
                  sig_34 <= sig_from_Fc;
               else
                  sig_34 <= sig_from_TmpA;
               end if;
               sig_to_Fd <= sig_34;
               if (sig_sel_TmpA = '0') then
                  sig_35 <= '1';
               else
                  sig_35 <= '0';
               end if;
               if (sig_35 = '1') then
                  sig_36 <= sig_from_Fd;
               else
                  sig_36 <= sig_from_TmpB;
               end if;
               sig_to_TmpA <= sig_36;
               if (sig_sel_TmpB = '0') then
                  sig_37 <= '1';
               else
                  sig_37 <= '0';
               end if;
               if (sig_37 = '1') then
                  sig_38 <= sig_from_TmpA;
               else
                  sig_38 <= sig_from_Xv;
               end if;
               sig_to_TmpB <= sig_38;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_39)) then
                  sig_40 <= '1';
               else
                  sig_40 <= '0';
               end if;
               if (unsigned(sig_sel_ToMALU) = unsigned(sig_41)) then
                  sig_42 <= '1';
               else
                  sig_42 <= '0';
               end if;
               if (sig_42 = '1') then
                  sig_43 <= sig_MALU_result;
               else
                  sig_43 <= sig_from_ToMALUShift;
               end if;
               if (sig_40 = '1') then
                  sig_44 <= sig_from_Xv;
               else
                  sig_44 <= sig_43;
               end if;
               sig_to_ToMALU <= sig_44;
               ready_int <= reg_ready;
               output_int <= sig_1;
               sig_en_out_Xv_int <= sig_en_Xv;
               sig_en_out_Yv_int <= sig_en_Yv;
               sig_en_out_Xp_int <= sig_en_Xp;
               sig_en_out_Yp_int <= sig_en_Yp;
               sig_en_out_Xfa_int <= sig_en_Xfa;
               sig_en_out_Yfa_int <= sig_en_Yfa;
               sig_en_out_Ga_int <= sig_en_Ga;
               sig_en_out_Gb_int <= sig_en_Gb;
               sig_en_out_Fa_int <= sig_en_Fa;
               sig_en_out_Fb_int <= sig_en_Fb;
               sig_en_out_Fc_int <= sig_en_Fc;
               sig_en_out_Fd_int <= sig_en_Fd;
               sig_en_out_TmpA_int <= sig_en_TmpA;
               sig_en_out_TmpB_int <= sig_en_TmpB;
               sig_en_out_ToMALU_int <= sig_en_ToMALU;
               reg_start_wire <= start_in;
               reg_next_wire <= next_in;
               reg_MALU_ready_wire <= sig_MALU_ready;
               sig_MALU_start <= '1';
               sig_MALU_mode <= '1';
               sig_MALU_plus_one <= '0';
               sig_sel_ToMALU <= sig_49;
               sig_en_ToMALU <= '1';
               reg_ToMALU_wire <= sig_to_ToMALU;
               sig_sel_Xv <= sig_54;
               sig_en_Xv <= '1';
               reg_Xv_wire <= sig_to_Xv;
               sig_sel_Yv <= '1';
               sig_en_Yv <= '1';
               reg_Yv_wire <= sig_to_Yv;
               sig_en_Xp <= '0';
               sig_sel_Xp <= '0';
               sig_en_Yp <= '0';
               sig_sel_Yp <= '0';
               sig_en_Xfa <= '0';
               sig_sel_Xfa <= '0';
               sig_en_Yfa <= '0';
               sig_sel_Yfa <= '0';
               sig_en_Ga <= '0';
               sig_sel_Ga <= '0';
               sig_en_Gb <= '0';
               sig_sel_Gb <= '0';
               sig_en_Fa <= '0';
               sig_sel_Fa <= '0';
               sig_en_Fb <= '0';
               sig_sel_Fb <= '0';
               sig_en_Fc <= '0';
               sig_sel_Fc <= '0';
               sig_en_Fd <= '0';
               sig_sel_Fd <= '0';
               sig_en_TmpA <= '0';
               sig_sel_TmpA <= '0';
               sig_sel_TmpB <= '1';
               sig_en_TmpB <= '1';
               reg_TmpB_wire <= sig_to_TmpB;
            when others=>
         end case;
      end process dpCMB;


   --controller reg
   fsmREG: process (CLK,RST)
      begin
         if (RST = '1') then
            STATE <= init1;
         elsif CLK' event and CLK = '1' then
            STATE <= STATE;
            case STATE is
               when init1 => 
                  if (sig_78 = '1') then
                          STATE <= init2;
                  else
                          STATE <= init1;
                  end if;
               when init2 => 
                  if (sig_79 = '1') then
                          STATE <= init2;
                  else
                     if (sig_80 = '1') then
                             STATE <= init3;
                     else
                             STATE <= init2;
                     end if;
                  end if;
               when init3 => 
                  if (sig_81 = '1') then
                          STATE <= init2;
                  else
                     if (sig_82 = '1') then
                             STATE <= init4;
                     else
                             STATE <= init3;
                     end if;
                  end if;
               when init4 => 
                  if (sig_83 = '1') then
                          STATE <= init2;
                  else
                     if (sig_84 = '1') then
                             STATE <= start;
                     else
                             STATE <= init4;
                     end if;
                  end if;
               when start => 
                       STATE <= distort1;
               when distort1 => 
                       STATE <= distort2;
               when distort2 => 
                       STATE <= distort3;
               when distort3 => 
                       STATE <= distort4;
               when distort4 => 
                       STATE <= distort5;
               when distort5 => 
                       STATE <= distort6;
               when distort6 => 
                       STATE <= distort7;
               when distort7 => 
                       STATE <= distort8;
               when distort8 => 
                       STATE <= miller_init1;
               when miller_init1 => 
                       STATE <= miller_init2;
               when miller_init2 => 
                       STATE <= startloop1;
               when startloop1 => 
                  if (sig_87 = '1') then
                          STATE <= finalexp1;
                  else
                     if (sig_88 = '1') then
                             STATE <= alambda1;
                     else
                             STATE <= dlambda1;
                     end if;
                  end if;
               when ready1 => 
                       STATE <= ready2;
               when ready2 => 
                  if (sig_85 = '1') then
                          STATE <= init2;
                  else
                     if (sig_86 = '1') then
                             STATE <= init1;
                     else
                             STATE <= ready2;
                     end if;
                  end if;
               when dlambda1 => 
                       STATE <= dlambda2;
               when dlambda2 => 
                       STATE <= dlambda3;
               when dlambda3 => 
                  if (sig_89 = '1') then
                          STATE <= dlambda3;
                  else
                          STATE <= coord1;
                  end if;
               when dlambda4 => 
                  if (sig_90 = '1') then
                          STATE <= coord1;
                  else
                          STATE <= coord1;
                  end if;
               when s => 
               when alambda1 => 
                       STATE <= alambda2;
               when alambda2 => 
                       STATE <= alambda3;
               when alambda3 => 
                       STATE <= alambda4;
               when alambda4 => 
                       STATE <= alambda5;
               when alambda5 => 
                       STATE <= alambda6;
               when alambda6 => 
                       STATE <= inv1;
               when alambda7 => 
                       STATE <= alambda8;
               when alambda8 => 
                       STATE <= alambda9;
               when alambda9 => 
                       STATE <= alambda10;
               when alambda10 => 
                       STATE <= alambda11;
               when alambda11 => 
                       STATE <= alambda12;
               when alambda12 => 
                       STATE <= alambda13;
               when alambda13 => 
                  if (sig_91 = '1') then
                          STATE <= alambda13;
                  else
                          STATE <= alambda14;
                  end if;
               when alambda14 => 
                       STATE <= alambda15;
               when alambda15 => 
                       STATE <= alambda16;
               when alambda16 => 
                       STATE <= alambda17;
               when alambda17 => 
                       STATE <= coord1;
               when inv1 => 
                       STATE <= inv2;
               when inv2 => 
                       STATE <= inv3;
               when inv3 => 
                       STATE <= inv4;
               when inv4 => 
                  if (sig_92 = '1') then
                          STATE <= inv4;
                  else
                          STATE <= inv5;
                  end if;
               when inv5 => 
                       STATE <= inv6;
               when inv6 => 
                  if (sig_93 = '1') then
                          STATE <= inv6;
                  else
                          STATE <= inv7;
                  end if;
               when inv7 => 
                       STATE <= inv8;
               when inv8 => 
                  if (sig_94 = '1') then
                          STATE <= inv8;
                  else
                          STATE <= inv9;
                  end if;
               when inv9 => 
                       STATE <= inv10;
               when inv10 => 
                  if (sig_95 = '1') then
                          STATE <= inv10;
                  else
                          STATE <= inv11;
                  end if;
               when inv11 => 
                       STATE <= inv12;
               when inv12 => 
                  if (sig_96 = '1') then
                          STATE <= inv12;
                  else
                          STATE <= inv13;
                  end if;
               when inv13 => 
                       STATE <= inv14;
               when inv14 => 
                  if (sig_97 = '1') then
                          STATE <= inv14;
                  else
                          STATE <= inv15;
                  end if;
               when inv15 => 
                       STATE <= inv16;
               when inv16 => 
                  if (sig_98 = '1') then
                          STATE <= inv16;
                  else
                          STATE <= inv17;
                  end if;
               when inv17 => 
                       STATE <= inv18;
               when inv18 => 
                       STATE <= inv19;
               when inv19 => 
                  if (sig_99 = '1') then
                          STATE <= inv21;
                  else
                          STATE <= inv20;
                  end if;
               when inv20 => 
                  if (sig_100 = '1') then
                          STATE <= inv20;
                  else
                          STATE <= inv19;
                  end if;
               when inv21 => 
                       STATE <= inv22;
               when inv22 => 
                  if (sig_101 = '1') then
                          STATE <= inv22;
                  else
                          STATE <= inv23;
                  end if;
               when inv23 => 
                       STATE <= inv24;
               when inv24 => 
                       STATE <= inv25;
               when inv25 => 
                  if (sig_102 = '1') then
                          STATE <= inv27;
                  else
                          STATE <= inv26;
                  end if;
               when inv26 => 
                  if (sig_103 = '1') then
                          STATE <= inv26;
                  else
                          STATE <= inv25;
                  end if;
               when inv27 => 
                       STATE <= inv28;
               when inv28 => 
                  if (sig_104 = '1') then
                          STATE <= inv28;
                  else
                          STATE <= inv29;
                  end if;
               when inv29 => 
                       STATE <= inv30;
               when inv30 => 
                       STATE <= inv31;
               when inv31 => 
                  if (sig_105 = '1') then
                          STATE <= inv33;
                  else
                          STATE <= inv32;
                  end if;
               when inv32 => 
                  if (sig_106 = '1') then
                          STATE <= inv32;
                  else
                          STATE <= inv31;
                  end if;
               when inv33 => 
                       STATE <= inv34;
               when inv34 => 
                  if (sig_107 = '1') then
                          STATE <= inv34;
                  else
                          STATE <= inv35;
                  end if;
               when inv35 => 
                       STATE <= inv36;
               when inv36 => 
                       STATE <= inv37;
               when inv37 => 
                  if (sig_108 = '1') then
                          STATE <= inv39;
                  else
                          STATE <= inv38;
                  end if;
               when inv38 => 
                  if (sig_109 = '1') then
                          STATE <= inv38;
                  else
                          STATE <= inv37;
                  end if;
               when inv39 => 
                       STATE <= inv40;
               when inv40 => 
                  if (sig_110 = '1') then
                          STATE <= inv40;
                  else
                          STATE <= inv41;
                  end if;
               when inv41 => 
                       STATE <= inv42;
               when inv42 => 
                  if (sig_111 = '1') then
                          STATE <= inv42;
                  else
                          STATE <= inv43;
                  end if;
               when inv43 => 
                       STATE <= inv44;
               when inv44 => 
                  if (sig_112 = '1') then
                          STATE <= inv44;
                  else
                          STATE <= inv45;
                  end if;
               when inv45 => 
                       STATE <= inv46;
               when inv46 => 
                       STATE <= inv47;
               when inv47 => 
                  if (sig_113 = '1') then
                          STATE <= inv49;
                  else
                          STATE <= inv48;
                  end if;
               when inv48 => 
                  if (sig_114 = '1') then
                          STATE <= inv48;
                  else
                          STATE <= inv47;
                  end if;
               when inv49 => 
                       STATE <= inv50;
               when inv50 => 
                  if (sig_115 = '1') then
                          STATE <= inv50;
                  else
                          STATE <= inv51;
                  end if;
               when inv51 => 
                       STATE <= inv52;
               when inv52 => 
                  if (sig_116 = '1') then
                          STATE <= inv52;
                  else
                          STATE <= inv53;
                  end if;
               when inv53 => 
                       STATE <= inv54;
               when inv54 => 
                  if (sig_117 = '1') then
                          STATE <= f2minv14;
                  else
                          STATE <= alambda7;
                  end if;
               when coord1 => 
                       STATE <= coord2;
               when coord2 => 
                  if (sig_118 = '1') then
                          STATE <= coord2;
                  else
                          STATE <= coord3;
                  end if;
               when coord3 => 
                  if (sig_119 = '1') then
                          STATE <= coord7;
                  else
                          STATE <= coord4;
                  end if;
               when coord4 => 
                       STATE <= coord5;
               when coord5 => 
                       STATE <= coord6;
               when coord6 => 
                       STATE <= coord7;
               when coord7 => 
                       STATE <= coord8;
               when coord8 => 
                       STATE <= coord9;
               when coord9 => 
                       STATE <= coord10;
               when coord10 => 
                       STATE <= coord11;
               when coord11 => 
                  if (sig_120 = '1') then
                          STATE <= coord11;
                  else
                          STATE <= coord12;
                  end if;
               when coord12 => 
                       STATE <= coord13;
               when coord13 => 
                       STATE <= coord14;
               when coord14 => 
                       STATE <= coord15;
               when coord15 => 
                       STATE <= coord16;
               when coord16 => 
                       STATE <= coord17;
               when coord17 => 
                       STATE <= coord18;
               when coord18 => 
                       STATE <= coord19;
               when coord19 => 
                  if (sig_121 = '1') then
                          STATE <= coord19;
                  else
                          STATE <= coord20;
                  end if;
               when coord20 => 
                       STATE <= coord21;
               when coord21 => 
                       STATE <= coord22;
               when coord22 => 
                       STATE <= coord23;
               when coord23 => 
                       STATE <= coord24;
               when coord24 => 
                       STATE <= coord25;
               when coord25 => 
                       STATE <= coord26;
               when coord26 => 
                       STATE <= coord27;
               when coord27 => 
                       STATE <= coord28;
               when coord28 => 
                       STATE <= coord29;
               when coord29 => 
                       STATE <= coord30;
               when coord30 => 
                       STATE <= coord31;
               when coord31 => 
                       STATE <= coord32;
               when coord32 => 
                       STATE <= coord33;
               when coord33 => 
                       STATE <= coord34;
               when coord34 => 
                       STATE <= coord35;
               when coord35 => 
                       STATE <= updatef1;
               when updatef1 => 
                  if (sig_122 = '1') then
                          STATE <= fsqrt1;
                  else
                          STATE <= fg1;
                  end if;
               when fsqrt1 => 
                       STATE <= fsqrt2;
               when fsqrt2 => 
                       STATE <= fsqrt3;
               when fsqrt3 => 
                       STATE <= fsqrt4;
               when fsqrt4 => 
                       STATE <= fsqrt5;
               when fsqrt5 => 
                       STATE <= fsqrt6;
               when fsqrt6 => 
                       STATE <= fsqrt7;
               when fsqrt7 => 
                       STATE <= fsqrt8;
               when fsqrt8 => 
                  if (sig_123 = '1') then
                          STATE <= fsqrt8;
                  else
                          STATE <= fsqrt9;
                  end if;
               when fsqrt9 => 
                       STATE <= fsqrt10;
               when fsqrt10 => 
                       STATE <= fsqrt11;
               when fsqrt11 => 
                       STATE <= fsqrt12;
               when fsqrt12 => 
                       STATE <= fsqrt13;
               when fsqrt13 => 
                       STATE <= fsqrt14;
               when fsqrt14 => 
                       STATE <= fsqrt15;
               when fsqrt15 => 
                  if (sig_124 = '1') then
                          STATE <= fsqrt15;
                  else
                          STATE <= fsqrt16;
                  end if;
               when fsqrt16 => 
                       STATE <= fsqrt17;
               when fsqrt17 => 
                       STATE <= fsqrt18;
               when fsqrt18 => 
                       STATE <= fsqrt19;
               when fsqrt19 => 
                       STATE <= fsqrt20;
               when fsqrt20 => 
                       STATE <= fsqrt21;
               when fsqrt21 => 
                       STATE <= fsqrt22;
               when fsqrt22 => 
                  if (sig_125 = '1') then
                          STATE <= fsqrt22;
                  else
                          STATE <= fsqrt23;
                  end if;
               when fsqrt23 => 
                       STATE <= fsqrt24;
               when fsqrt24 => 
                       STATE <= fsqrt25;
               when fsqrt25 => 
                       STATE <= fsqrt26;
               when fsqrt26 => 
                  if (sig_126 = '1') then
                          STATE <= fsqrt26;
                  else
                          STATE <= fsqrt27;
                  end if;
               when fsqrt27 => 
                       STATE <= fsqrt28;
               when fsqrt28 => 
                       STATE <= fsqrt29;
               when fsqrt29 => 
                       STATE <= fsqrt30;
               when fsqrt30 => 
                       STATE <= fsqrt31;
               when fsqrt31 => 
                       STATE <= fsqrt32;
               when fsqrt32 => 
                       STATE <= fg1;
               when fg1 => 
                       STATE <= fg2;
               when fg2 => 
                       STATE <= fg3;
               when fg3 => 
                       STATE <= fg4;
               when fg4 => 
                       STATE <= fg5;
               when fg5 => 
                       STATE <= fg6;
               when fg6 => 
                       STATE <= fg7;
               when fg7 => 
                  if (sig_127 = '1') then
                          STATE <= fg7;
                  else
                          STATE <= fg8;
                  end if;
               when fg8 => 
                       STATE <= fg9;
               when fg9 => 
                       STATE <= fg10;
               when fg10 => 
                       STATE <= fg11;
               when fg11 => 
                       STATE <= fg12;
               when fg12 => 
                       STATE <= fg13;
               when fg13 => 
                       STATE <= fg14;
               when fg14 => 
                       STATE <= fg15;
               when fg15 => 
                       STATE <= fg16;
               when fg16 => 
                       STATE <= fg17;
               when fg17 => 
                       STATE <= fg18;
               when fg18 => 
                       STATE <= fg19;
               when fg19 => 
                       STATE <= fg20;
               when fg20 => 
                       STATE <= fg21;
               when fg21 => 
                       STATE <= fg22;
               when fg22 => 
                       STATE <= fg23;
               when fg23 => 
                  if (sig_128 = '1') then
                          STATE <= fg23;
                  else
                          STATE <= fg24;
                  end if;
               when fg24 => 
                       STATE <= fg25;
               when fg25 => 
                       STATE <= fg26;
               when fg26 => 
                       STATE <= fg27;
               when fg27 => 
                       STATE <= fg28;
               when fg28 => 
                       STATE <= fg29;
               when fg29 => 
                       STATE <= fg30;
               when fg30 => 
                  if (sig_129 = '1') then
                          STATE <= fg30;
                  else
                          STATE <= fg31;
                  end if;
               when fg31 => 
                       STATE <= fg32;
               when fg32 => 
                       STATE <= fg33;
               when fg33 => 
                       STATE <= fg34;
               when fg34 => 
                       STATE <= fg35;
               when fg35 => 
                  if (sig_130 = '1') then
                          STATE <= fg35;
                  else
                          STATE <= fg36;
                  end if;
               when fg36 => 
                       STATE <= fg37;
               when fg37 => 
                       STATE <= fg38;
               when fg38 => 
                       STATE <= fg39;
               when fg39 => 
                       STATE <= fg40;
               when fg40 => 
                       STATE <= fg41;
               when fg41 => 
                       STATE <= fg42;
               when fg42 => 
                       STATE <= fg43;
               when fg43 => 
                       STATE <= fg44;
               when fg44 => 
                       STATE <= fg45;
               when fg45 => 
                       STATE <= fg46;
               when fg46 => 
                  if (sig_131 = '1') then
                          STATE <= fg46;
                  else
                          STATE <= fg47;
                  end if;
               when fg47 => 
                       STATE <= fg48;
               when fg48 => 
                       STATE <= fg49;
               when fg49 => 
                       STATE <= fg50;
               when fg50 => 
                       STATE <= fg51;
               when fg51 => 
                       STATE <= fg52;
               when fg52 => 
                       STATE <= fg53;
               when fg53 => 
                       STATE <= fg54;
               when fg54 => 
                       STATE <= fg55;
               when fg55 => 
                       STATE <= fg56;
               when fg56 => 
                       STATE <= fg57;
               when fg57 => 
                       STATE <= fg58;
               when fg58 => 
                       STATE <= fg59;
               when fg59 => 
                  if (sig_132 = '1') then
                          STATE <= fg59;
                  else
                          STATE <= fg60;
                  end if;
               when fg60 => 
                       STATE <= fg61;
               when fg61 => 
                       STATE <= fg62;
               when fg62 => 
                       STATE <= fg63;
               when fg63 => 
                       STATE <= fg64;
               when fg64 => 
                       STATE <= fg65;
               when fg65 => 
                       STATE <= fg66;
               when fg66 => 
                       STATE <= fg67;
               when fg67 => 
                  if (sig_135 = '1') then
                          STATE <= startloop1;
                  else
                          STATE <= startloop1;
                  end if;
               when finalexp1 => 
                       STATE <= finalexp2;
               when finalexp2 => 
                       STATE <= finalexp3;
               when finalexp3 => 
                       STATE <= finalexp4;
               when finalexp4 => 
                       STATE <= finalexp5;
               when finalexp5 => 
                  if (sig_136 = '1') then
                          STATE <= finalexp5;
                  else
                          STATE <= finalexp6;
                  end if;
               when finalexp6 => 
                       STATE <= finalexp7;
               when finalexp7 => 
                       STATE <= finalexp8;
               when finalexp8 => 
                       STATE <= finalexp9;
               when finalexp9 => 
                  if (sig_137 = '1') then
                          STATE <= finalexp9;
                  else
                          STATE <= finalexp10;
                  end if;
               when finalexp10 => 
                       STATE <= finalexp11;
               when finalexp11 => 
                       STATE <= finalexp12;
               when finalexp12 => 
                       STATE <= finalexp13;
               when finalexp13 => 
                  if (sig_138 = '1') then
                          STATE <= finalexp13;
                  else
                          STATE <= finalexp14;
                  end if;
               when finalexp14 => 
                       STATE <= finalexp15;
               when finalexp15 => 
                       STATE <= finalexp16;
               when finalexp16 => 
                       STATE <= finalexp17;
               when finalexp17 => 
                  if (sig_139 = '1') then
                          STATE <= finalexp17;
                  else
                          STATE <= finalexp18;
                  end if;
               when finalexp18 => 
                       STATE <= finalexp19;
               when finalexp19 => 
                       STATE <= finalexp20;
               when finalexp20 => 
                       STATE <= finalexp21;
               when finalexp21 => 
                       STATE <= finalexp22;
               when finalexp22 => 
                       STATE <= finalexp23;
               when finalexp23 => 
                       STATE <= finalexp24;
               when finalexp24 => 
                       STATE <= finalexp25;
               when finalexp25 => 
                       STATE <= finalexp26;
               when finalexp26 => 
                       STATE <= finalexp27;
               when finalexp27 => 
                       STATE <= finalexp28;
               when finalexp28 => 
                       STATE <= finalexp29;
               when finalexp29 => 
                       STATE <= finalexp30;
               when finalexp30 => 
                       STATE <= finalexp31;
               when finalexp31 => 
                       STATE <= finalexp32;
               when finalexp32 => 
                       STATE <= finalexp33;
               when finalexp33 => 
                       STATE <= finalexp34;
               when finalexp34 => 
                       STATE <= finalexp35;
               when finalexp35 => 
                       STATE <= finalexp36;
               when finalexp36 => 
                       STATE <= finalexp37;
               when finalexp37 => 
                       STATE <= finalexp38;
               when finalexp38 => 
                       STATE <= finalexp39;
               when finalexp39 => 
                       STATE <= finalexp40;
               when finalexp40 => 
                       STATE <= finalexp41;
               when finalexp41 => 
                  if (sig_140 = '1') then
                          STATE <= finalexp41;
                  else
                          STATE <= finalexp42;
                  end if;
               when finalexp42 => 
                       STATE <= finalexp43;
               when finalexp43 => 
                       STATE <= finalexp44;
               when finalexp44 => 
                       STATE <= finalexp45;
               when finalexp45 => 
                       STATE <= finalexp46;
               when finalexp46 => 
                  if (sig_141 = '1') then
                          STATE <= finalexp46;
                  else
                          STATE <= finalexp47;
                  end if;
               when finalexp47 => 
                       STATE <= finalexp48;
               when finalexp48 => 
                       STATE <= finalexp49;
               when finalexp49 => 
                       STATE <= finalexp50;
               when finalexp50 => 
                       STATE <= finalexp51;
               when finalexp51 => 
                  if (sig_142 = '1') then
                          STATE <= finalexp51;
                  else
                          STATE <= finalexp52;
                  end if;
               when finalexp52 => 
                       STATE <= finalexp53;
               when finalexp53 => 
                       STATE <= finalexp54;
               when finalexp54 => 
                       STATE <= finalexp55;
               when finalexp55 => 
                       STATE <= finalexp56;
               when finalexp56 => 
                       STATE <= finalexp57;
               when finalexp57 => 
                       STATE <= finalexp58;
               when finalexp58 => 
                       STATE <= finalexp59;
               when finalexp59 => 
                       STATE <= finalexp60;
               when finalexp60 => 
                       STATE <= finalexp61;
               when finalexp61 => 
                       STATE <= finalexp62;
               when finalexp62 => 
                       STATE <= finalexp63;
               when finalexp63 => 
                       STATE <= f2minv1;
               when finalexp64 => 
                       STATE <= finalexp65;
               when finalexp65 => 
                       STATE <= finalexp66;
               when finalexp66 => 
                       STATE <= finalexp67;
               when finalexp67 => 
                       STATE <= finalexp68;
               when finalexp68 => 
                       STATE <= finalexp69;
               when finalexp69 => 
                       STATE <= finalexp70;
               when finalexp70 => 
                       STATE <= finalexp71;
               when finalexp71 => 
                       STATE <= finalexp72;
               when finalexp72 => 
                       STATE <= finalexp73;
               when finalexp73 => 
                       STATE <= finalexp74;
               when finalexp74 => 
                       STATE <= finalexp75;
               when finalexp75 => 
                       STATE <= finalexp76;
               when finalexp76 => 
                       STATE <= finalexp77;
               when finalexp77 => 
                       STATE <= finalexp78;
               when finalexp78 => 
                       STATE <= finalexp79;
               when finalexp79 => 
                       STATE <= finalexp80;
               when finalexp80 => 
                       STATE <= f2mmult1;
               when f4mpow1 => 
                       STATE <= f4mpow2;
               when f4mpow2 => 
                       STATE <= f4mpow3;
               when f4mpow3 => 
                       STATE <= f4mpow4;
               when f4mpow4 => 
                       STATE <= f4mpow5;
               when f4mpow5 => 
                       STATE <= f4mpow6;
               when f4mpow6 => 
                       STATE <= f4mpow7;
               when f4mpow7 => 
                       STATE <= f4mpow8;
               when f4mpow8 => 
                       STATE <= f4mpow9;
               when f4mpow9 => 
                       STATE <= f4mpow10;
               when f4mpow10 => 
                       STATE <= f4mpow11;
               when f4mpow11 => 
                       STATE <= f4mpow12;
               when f4mpow12 => 
                       STATE <= f4mpow13;
               when f4mpow13 => 
                       STATE <= f4mpow14;
               when f4mpow14 => 
                       STATE <= f4mpow15;
               when f4mpow15 => 
                  if (sig_143 = '1') then
                          STATE <= f4mpow15;
                  else
                          STATE <= f4mpow16;
                  end if;
               when f4mpow16 => 
                       STATE <= f4mpow17;
               when f4mpow17 => 
                       STATE <= f4mpow18;
               when f4mpow18 => 
                       STATE <= f4mpow19;
               when f4mpow19 => 
                       STATE <= f4mpow20;
               when f4mpow20 => 
                       STATE <= f4mpow21;
               when f4mpow21 => 
                  if (sig_144 = '1') then
                          STATE <= f4mpow21;
                  else
                          STATE <= f4mpow22;
                  end if;
               when f4mpow22 => 
                       STATE <= f4mpow23;
               when f4mpow23 => 
                       STATE <= f4mpow24;
               when f4mpow24 => 
                  if (sig_145 = '1') then
                          STATE <= f4mpow24;
                  else
                          STATE <= f4mpow25;
                  end if;
               when f4mpow25 => 
                       STATE <= f4mpow26;
               when f4mpow26 => 
                       STATE <= f4mpow27;
               when f4mpow27 => 
                       STATE <= f4mpow28;
               when f4mpow28 => 
                  if (sig_146 = '1') then
                          STATE <= f4mpow28;
                  else
                          STATE <= f4mpow29;
                  end if;
               when f4mpow29 => 
                       STATE <= f4mpow30;
               when f4mpow30 => 
                       STATE <= f4mpow31;
               when f4mpow31 => 
                       STATE <= f4mpow32;
               when f4mpow32 => 
                       STATE <= f4mpow33;
               when f4mpow33 => 
                       STATE <= f4mpow34;
               when f4mpow34 => 
                  if (sig_147 = '1') then
                          STATE <= f4mpow34;
                  else
                          STATE <= f4mpow35;
                  end if;
               when f4mpow35 => 
                       STATE <= f4mpow36;
               when f4mpow36 => 
                       STATE <= f4mpow37;
               when f4mpow37 => 
                  if (sig_148 = '1') then
                          STATE <= f4mpow37;
                  else
                          STATE <= f4mpow38;
                  end if;
               when f4mpow38 => 
                       STATE <= f4mpow39;
               when f4mpow39 => 
                       STATE <= f4mpow40;
               when f4mpow40 => 
                  if (sig_149 = '1') then
                          STATE <= f4mpow40;
                  else
                          STATE <= f4mpow41;
                  end if;
               when f4mpow41 => 
                       STATE <= f4mpow42;
               when f4mpow42 => 
                       STATE <= f4mpow43;
               when f4mpow43 => 
                       STATE <= f4mpow44;
               when f4mpow44 => 
                       STATE <= f4mpow45;
               when f4mpow45 => 
                       STATE <= f4mpow46;
               when f4mpow46 => 
                       STATE <= f4mpow47fix;
               when f4mpow47 => 
                       STATE <= f4mpow48;
               when f4mpow48 => 
                       STATE <= f4mpow49;
               when f4mpow49 => 
                       STATE <= f4mpow50;
               when f4mpow50 => 
                       STATE <= f4mpow51;
               when f4mpow51 => 
                       STATE <= f4mpow52;
               when f4mpow52 => 
                       STATE <= f4mpow53;
               when f4mpow53 => 
                       STATE <= f4mpow54;
               when f4mpow54 => 
                       STATE <= f4mpow55;
               when f4mpow55 => 
                       STATE <= f4mpow56;
               when f4mpow56 => 
                       STATE <= f4mpow57;
               when f4mpow57 => 
                       STATE <= f4mpow58;
               when f4mpow58 => 
                       STATE <= f4mpow59;
               when f4mpow59 => 
                       STATE <= f4mpow60;
               when f4mpow60 => 
                       STATE <= f4mpow61;
               when f4mpow61 => 
                       STATE <= f4mpow62;
               when f4mpow62 => 
                       STATE <= f4msqrt1;
               when f4mpow47fix => 
                       STATE <= f4mpow47;
               when f4msqrt1 => 
                       STATE <= f4msqrt2;
               when f4msqrt2 => 
                  if (sig_150 = '1') then
                          STATE <= f4mmult1;
                  else
                          STATE <= f4msqrt3;
                  end if;
               when f4msqrt3 => 
                       STATE <= f4msqrt4;
               when f4msqrt4 => 
                       STATE <= f4msqrt5;
               when f4msqrt5 => 
                  if (sig_151 = '1') then
                          STATE <= f4msqrt5;
                  else
                          STATE <= f4msqrt6;
                  end if;
               when f4msqrt6 => 
                       STATE <= f4msqrt7;
               when f4msqrt7 => 
                       STATE <= f4msqrt8;
               when f4msqrt8 => 
                  if (sig_152 = '1') then
                          STATE <= f4msqrt8;
                  else
                          STATE <= f4msqrt9;
                  end if;
               when f4msqrt9 => 
                       STATE <= f4msqrt10;
               when f4msqrt10 => 
                       STATE <= f4msqrt11;
               when f4msqrt11 => 
                  if (sig_153 = '1') then
                          STATE <= f4msqrt11;
                  else
                          STATE <= f4msqrt12;
                  end if;
               when f4msqrt12 => 
                       STATE <= f4msqrt13;
               when f4msqrt13 => 
                       STATE <= f4msqrt14;
               when f4msqrt14 => 
                  if (sig_154 = '1') then
                          STATE <= f4msqrt14;
                  else
                          STATE <= f4msqrt15;
                  end if;
               when f4msqrt15 => 
                       STATE <= f4msqrt16;
               when f4msqrt16 => 
                       STATE <= f4msqrt17;
               when f4msqrt17 => 
                       STATE <= f4msqrt18;
               when f4msqrt18 => 
                       STATE <= f4msqrt19;
               when f4msqrt19 => 
                       STATE <= f4msqrt20;
               when f4msqrt20 => 
                       STATE <= f4msqrt21;
               when f4msqrt21 => 
                       STATE <= f4msqrt22;
               when f4msqrt22 => 
                       STATE <= f4msqrt23;
               when f4msqrt23 => 
                       STATE <= f4msqrt24;
               when f4msqrt24 => 
                       STATE <= f4msqrt25;
               when f4msqrt25 => 
                       STATE <= f4msqrt26;
               when f4msqrt26 => 
                       STATE <= f4msqrt27fix;
               when f4msqrt27 => 
                       STATE <= f4msqrt28;
               when f4msqrt28 => 
                       STATE <= f4msqrt29;
               when f4msqrt29 => 
                       STATE <= f4msqrt30;
               when f4msqrt30 => 
                       STATE <= f4msqrt31;
               when f4msqrt31 => 
                       STATE <= f4msqrt32;
               when f4msqrt32 => 
                       STATE <= f4msqrt2;
               when f4msqrt27fix => 
                       STATE <= f4msqrt27;
               when f4mmult1 => 
                       STATE <= f4mmult2;
               when f4mmult2 => 
                       STATE <= f4mmult3;
               when f4mmult3 => 
                       STATE <= f4mmult4;
               when f4mmult4 => 
                       STATE <= f4mmult5;
               when f4mmult5 => 
                       STATE <= f4mmult6;
               when f4mmult6 => 
                       STATE <= f4mmult7;
               when f4mmult7 => 
                       STATE <= f4mmult8;
               when f4mmult8 => 
                       STATE <= f4mmult9;
               when f4mmult9 => 
                       STATE <= f4mmult10;
               when f4mmult10 => 
                  if (sig_155 = '1') then
                          STATE <= f4mmult10;
                  else
                          STATE <= f4mmult11;
                  end if;
               when f4mmult11 => 
                       STATE <= f4mmult12;
               when f4mmult12 => 
                       STATE <= f4mmult13;
               when f4mmult13 => 
                       STATE <= f4mmult14;
               when f4mmult14 => 
                       STATE <= f4mmult15;
               when f4mmult15 => 
                       STATE <= f4mmult16;
               when f4mmult16 => 
                       STATE <= f4mmult17;
               when f4mmult17 => 
                       STATE <= f4mmult18;
               when f4mmult18 => 
                       STATE <= f4mmult19;
               when f4mmult19 => 
                  if (sig_156 = '1') then
                          STATE <= f4mmult19;
                  else
                          STATE <= f4mmult20;
                  end if;
               when f4mmult20 => 
                       STATE <= f4mmult21;
               when f4mmult21 => 
                       STATE <= f4mmult22;
               when f4mmult22 => 
                       STATE <= f4mmult23;
               when f4mmult23 => 
                       STATE <= f4mmult24;
               when f4mmult24 => 
                       STATE <= f4mmult25;
               when f4mmult25 => 
                       STATE <= f4mmult26;
               when f4mmult26 => 
                       STATE <= f4mmult27;
               when f4mmult27 => 
                       STATE <= f4mmult28;
               when f4mmult28 => 
                       STATE <= f4mmult29;
               when f4mmult29 => 
                       STATE <= f4mmult30;
               when f4mmult30 => 
                       STATE <= f4mmult31;
               when f4mmult31 => 
                       STATE <= f4mmult32;
               when f4mmult32 => 
                       STATE <= f4mmult33;
               when f4mmult33 => 
                       STATE <= f4mmult34;
               when f4mmult34 => 
                       STATE <= f4mmult35;
               when f4mmult35 => 
                       STATE <= f4mmult36;
               when f4mmult36 => 
                  if (sig_157 = '1') then
                          STATE <= f4mmult36;
                  else
                          STATE <= f4mmult37;
                  end if;
               when f4mmult37 => 
                       STATE <= f4mmult38;
               when f4mmult38 => 
                       STATE <= f4mmult39;
               when f4mmult39 => 
                       STATE <= f4mmult40;
               when f4mmult40 => 
                  if (sig_158 = '1') then
                          STATE <= f4mmult40;
                  else
                          STATE <= f4mmult41;
                  end if;
               when f4mmult41 => 
                       STATE <= f4mmult42;
               when f4mmult42 => 
                       STATE <= f4mmult43;
               when f4mmult43 => 
                       STATE <= f4mmult44;
               when f4mmult44 => 
                       STATE <= f4mmult45;
               when f4mmult45 => 
                  if (sig_159 = '1') then
                          STATE <= f4mmult45;
                  else
                          STATE <= f4mmult46;
                  end if;
               when f4mmult46 => 
                       STATE <= f4mmult47;
               when f4mmult47 => 
                       STATE <= f4mmult48;
               when f4mmult48 => 
                  if (sig_160 = '1') then
                          STATE <= f4mmult48;
                  else
                          STATE <= f4mmult49;
                  end if;
               when f4mmult49 => 
                       STATE <= f4mmult50;
               when f4mmult50 => 
                       STATE <= f4mmult51;
               when f4mmult51 => 
                  if (sig_161 = '1') then
                          STATE <= f4mmult51;
                  else
                          STATE <= f4mmult52;
                  end if;
               when f4mmult52 => 
                       STATE <= f4mmult53;
               when f4mmult53 => 
                       STATE <= f4mmult54;
               when f4mmult54 => 
                       STATE <= f4mmult55;
               when f4mmult55 => 
                       STATE <= f4mmult56;
               when f4mmult56 => 
                       STATE <= f4mmult57;
               when f4mmult57 => 
                  if (sig_162 = '1') then
                          STATE <= f4mmult57;
                  else
                          STATE <= f4mmult58;
                  end if;
               when f4mmult58 => 
                       STATE <= f4mmult59;
               when f4mmult59 => 
                       STATE <= f4mmult60;
               when f4mmult60 => 
                       STATE <= f4mmult61;
               when f4mmult61 => 
                       STATE <= f4mmult62;
               when f4mmult62 => 
                  if (sig_163 = '1') then
                          STATE <= f4mmult62;
                  else
                          STATE <= f4mmult63;
                  end if;
               when f4mmult63 => 
                       STATE <= f4mmult64;
               when f4mmult64 => 
                       STATE <= f4mmult65;
               when f4mmult65 => 
                       STATE <= f4mmult66;
               when f4mmult66 => 
                       STATE <= f4mmult67;
               when f4mmult67 => 
                       STATE <= f4mmult68;
               when f4mmult68 => 
                       STATE <= f4mmult69;
               when f4mmult69 => 
                       STATE <= f4mmult70;
               when f4mmult70 => 
                       STATE <= f4mmult71;
               when f4mmult71 => 
                       STATE <= f4mmfix1;
               when f4mmult72 => 
               when f4mmult73 => 
                       STATE <= f4mmult74;
               when f4mmult74 => 
                       STATE <= f4mmfix4;
               when f4mmult75 => 
                       STATE <= f4mmult76;
               when f4mmult76 => 
                       STATE <= f4mmult77;
               when f4mmult77 => 
                       STATE <= f4mmult78;
               when f4mmult78 => 
                       STATE <= f4mmult79;
               when f4mmult79 => 
                       STATE <= f4mmult80;
               when f4mmult80 => 
                       STATE <= f4mmult81;
               when f4mmult81 => 
                       STATE <= f4mmult82;
               when f4mmult82 => 
                       STATE <= f4mmult83;
               when f4mmult83 => 
                       STATE <= f4mmult84;
               when f4mmult84 => 
                       STATE <= f4mmult85;
               when f4mmult85 => 
                       STATE <= f4mmult86;
               when f4mmult86 => 
                       STATE <= f4mmult87;
               when f4mmult87 => 
                       STATE <= f4mmult88;
               when f4mmult88 => 
                       STATE <= f4mmult89;
               when f4mmult89 => 
                       STATE <= f4mmult90;
               when f4mmult90 => 
                       STATE <= f4mmult91;
               when f4mmult91 => 
                       STATE <= f4mmult92;
               when f4mmult92 => 
                       STATE <= f4mmult93;
               when f4mmult93 => 
                       STATE <= f4mmult94;
               when f4mmult94 => 
                       STATE <= f4mmult95;
               when f4mmult95 => 
                       STATE <= f4mmult96;
               when f4mmult96 => 
                       STATE <= ready1;
               when f4mmfix1 => 
                       STATE <= f4mmfix2;
               when f4mmfix2 => 
                       STATE <= f4mmfix3;
               when f4mmfix3 => 
                       STATE <= f4mmult73;
               when f4mmfix4 => 
                       STATE <= f4mmfix5;
               when f4mmfix5 => 
                       STATE <= f4mmult75;
               when f2mmult1 => 
                       STATE <= f2mmult2;
               when f2mmult2 => 
                  if (sig_164 = '1') then
                          STATE <= f4mpow1;
                  else
                          STATE <= f2mmult3;
                  end if;
               when f2mmult3 => 
                       STATE <= f2mmult4;
               when f2mmult4 => 
                       STATE <= f2mmult5;
               when f2mmult5 => 
                       STATE <= f2mmult6;
               when f2mmult6 => 
                       STATE <= f2mmult7;
               when f2mmult7 => 
                       STATE <= f2mmult8;
               when f2mmult8 => 
                       STATE <= f2mmult9;
               when f2mmult9 => 
                  if (sig_165 = '1') then
                          STATE <= f2mmult9;
                  else
                          STATE <= f2mmult10;
                  end if;
               when f2mmult10 => 
                       STATE <= f2mmult11;
               when f2mmult11 => 
                       STATE <= f2mmult12;
               when f2mmult12 => 
                       STATE <= f2mmult13;
               when f2mmult13 => 
                       STATE <= f2mmult14;
               when f2mmult14 => 
                       STATE <= f2mmult15;
               when f2mmult15 => 
                       STATE <= f2mmult16;
               when f2mmult16 => 
                  if (sig_166 = '1') then
                          STATE <= f2mmult16;
                  else
                          STATE <= f2mmult17;
                  end if;
               when f2mmult17 => 
                       STATE <= f2mmult18;
               when f2mmult18 => 
                       STATE <= f2mmult19;
               when f2mmult19 => 
                  if (sig_167 = '1') then
                          STATE <= f2mmult19;
                  else
                          STATE <= f2mmult20;
                  end if;
               when f2mmult20 => 
                       STATE <= f2mmult21;
               when f2mmult21 => 
                       STATE <= f2mmult22;
               when f2mmult22 => 
                       STATE <= f2mmult23;
               when f2mmult23 => 
                       STATE <= f2mmult24;
               when f2mmult24 => 
                       STATE <= f2mmult25;
               when f2mmult25 => 
                       STATE <= f2mmult26;
               when f2mmult26 => 
                       STATE <= f2mmult27;
               when f2mmult27 => 
                       STATE <= f2mmult28;
               when f2mmult28 => 
                       STATE <= f2mmult29;
               when f2mmult29 => 
                       STATE <= f2mmult2;
               when f2minv1 => 
                       STATE <= f2minv2;
               when f2minv2 => 
                       STATE <= f2minv3;
               when f2minv3 => 
                       STATE <= f2minv4;
               when f2minv4 => 
                       STATE <= f2minv5;
               when f2minv5 => 
                       STATE <= f2minv6;
               when f2minv6 => 
                  if (sig_168 = '1') then
                          STATE <= f2minv6;
                  else
                          STATE <= f2minv7;
                  end if;
               when f2minv7 => 
                       STATE <= f2minv8;
               when f2minv8 => 
                       STATE <= f2minv9;
               when f2minv9 => 
                       STATE <= f2minv10;
               when f2minv10 => 
                  if (sig_169 = '1') then
                          STATE <= f2minv10;
                  else
                          STATE <= f2minv11;
                  end if;
               when f2minv11 => 
                       STATE <= f2minv12;
               when f2minv12 => 
                       STATE <= f2minv13;
               when f2minv13 => 
                       STATE <= inv1;
               when f2minv14 => 
                       STATE <= f2minv15;
               when f2minv15 => 
                  if (sig_170 = '1') then
                          STATE <= f2minv15;
                  else
                          STATE <= f2minv16;
                  end if;
               when f2minv16 => 
                       STATE <= f2minv17;
               when f2minv17 => 
                       STATE <= f2minv18;
               when f2minv18 => 
                  if (sig_171 = '1') then
                          STATE <= f2minv18;
                  else
                          STATE <= f2minv19;
                  end if;
               when f2minv19 => 
                       STATE <= finalexp64;
               when others=>
            end case;
         end if;
      end process fsmREG;


   --controller cmb
   fsmCMB: process (reg_Xv,reg_Yv,reg_Xp,reg_Yp,reg_Xfa,reg_Yfa,reg_Ga,reg_Gb,reg_Fa,reg_Fb
,reg_Fc,reg_Fd,reg_TmpA,reg_TmpB,reg_ToMALU,reg_MALU_ready,reg_counter_miller,reg_counter_misc,reg_add,reg_start
,reg_next,reg_ready,sig_MALU_A,sig_MALU_B,sig_MALU_start,sig_MALU_mode,sig_MALU_plus_one,sig_MALU_result,sig_MALU_ready,sig_en_Xv
,sig_en_Yv,sig_en_Xp,sig_en_Yp,sig_en_Xfa,sig_en_Yfa,sig_en_Ga,sig_en_Gb,sig_en_Fa,sig_en_Fb,sig_en_Fc
,sig_en_Fd,sig_en_TmpA,sig_en_TmpB,sig_en_ToMALU,sig_sel_Xv,sig_sel_Yv,sig_sel_Xp,sig_sel_Yp,sig_sel_Xfa,sig_sel_Yfa
,sig_sel_Ga,sig_sel_Gb,sig_sel_Fa,sig_sel_Fb,sig_sel_Fc,sig_sel_Fd,sig_sel_TmpA,sig_sel_TmpB,sig_sel_ToMALU,sig_to_Xv
,sig_to_Yv,sig_to_Xp,sig_to_Yp,sig_to_Xfa,sig_to_Yfa,sig_to_Ga,sig_to_Gb,sig_to_Fa,sig_to_Fb,sig_to_Fc
,sig_to_Fd,sig_to_TmpA,sig_to_TmpB,sig_to_ToMALU,sig_from_Xv,sig_from_Yv,sig_from_Xp,sig_from_Yp,sig_from_Xfa,sig_from_Yfa
,sig_from_Ga,sig_from_Gb,sig_from_Fa,sig_from_Fb,sig_from_Fc,sig_from_Fd,sig_from_TmpA,sig_from_TmpB,sig_from_ToMALU,sig_from_ToMALUShift
,sig_from_Input,sig_0,sig_1,sig_2,sig_3,sig_4,sig_6,sig_8,sig_10,sig_11
,sig_12,sig_13,sig_14,sig_15,sig_16,sig_17,sig_18,sig_19,sig_20,sig_21
,sig_22,sig_23,sig_24,sig_25,sig_26,sig_27,sig_28,sig_29,sig_30,sig_31
,sig_32,sig_33,sig_34,sig_35,sig_36,sig_37,sig_38,sig_40,sig_42,sig_43
,sig_44,sig_56,sig_57,sig_58,sig_59,sig_60,sig_61,sig_62,sig_64,sig_65
,sig_66,sig_67,sig_68,sig_69,sig_70,sig_71,sig_72,sig_73,sig_74,sig_75
,ready_int,output_int,sig_en_out_Xv_int,sig_en_out_Yv_int,sig_en_out_Xp_int,sig_en_out_Yp_int,sig_en_out_Xfa_int,sig_en_out_Yfa_int,sig_en_out_Ga_int,sig_en_out_Gb_int
,sig_en_out_Fa_int,sig_en_out_Fb_int,sig_en_out_Fc_int,sig_en_out_Fd_int,sig_en_out_TmpA_int,sig_en_out_TmpB_int,sig_en_out_ToMALU_int,sig_78,sig_79,sig_80
,sig_81,sig_82,sig_83,sig_84,sig_85,sig_86,sig_87,sig_88,sig_89,sig_90
,sig_91,sig_92,sig_93,sig_94,sig_95,sig_96,sig_97,sig_98,sig_99,sig_100
,sig_101,sig_102,sig_103,sig_104,sig_105,sig_106,sig_107,sig_108,sig_109,sig_110
,sig_111,sig_112,sig_113,sig_114,sig_115,sig_116,sig_117,sig_118,sig_119,sig_120
,sig_121,sig_122,sig_123,sig_124,sig_125,sig_126,sig_127,sig_128,sig_129,sig_130
,sig_131,sig_132,sig_133,sig_134,sig_135,sig_136,sig_137,sig_138,sig_139,sig_140
,sig_141,sig_142,sig_143,sig_144,sig_145,sig_146,sig_147,sig_148,sig_149,sig_150
,sig_151,sig_152,sig_153,sig_154,sig_155,sig_156,sig_157,sig_158,sig_159,sig_160
,sig_161,sig_162,sig_163,sig_164,sig_165,sig_166,sig_167,sig_168,sig_169,sig_170
,sig_171,input,start_in,next_in,cmd,STATE)
      begin
      sig_78 <= '0';
      sig_79 <= '0';
      sig_80 <= '0';
      sig_81 <= '0';
      sig_82 <= '0';
      sig_83 <= '0';
      sig_84 <= '0';
      sig_85 <= '0';
      sig_86 <= '0';
      sig_87 <= '0';
      sig_88 <= '0';
      sig_89 <= '0';
      sig_90 <= '0';
      sig_91 <= '0';
      sig_92 <= '0';
      sig_93 <= '0';
      sig_94 <= '0';
      sig_95 <= '0';
      sig_96 <= '0';
      sig_97 <= '0';
      sig_98 <= '0';
      sig_99 <= '0';
      sig_100 <= '0';
      sig_101 <= '0';
      sig_102 <= '0';
      sig_103 <= '0';
      sig_104 <= '0';
      sig_105 <= '0';
      sig_106 <= '0';
      sig_107 <= '0';
      sig_108 <= '0';
      sig_109 <= '0';
      sig_110 <= '0';
      sig_111 <= '0';
      sig_112 <= '0';
      sig_113 <= '0';
      sig_114 <= '0';
      sig_115 <= '0';
      sig_116 <= '0';
      sig_117 <= '0';
      sig_118 <= '0';
      sig_119 <= '0';
      sig_120 <= '0';
      sig_121 <= '0';
      sig_122 <= '0';
      sig_123 <= '0';
      sig_124 <= '0';
      sig_125 <= '0';
      sig_126 <= '0';
      sig_127 <= '0';
      sig_128 <= '0';
      sig_129 <= '0';
      sig_130 <= '0';
      sig_131 <= '0';
      sig_132 <= '0';
      sig_133 <= '0';
      sig_134 <= '0';
      sig_135 <= '0';
      sig_136 <= '0';
      sig_137 <= '0';
      sig_138 <= '0';
      sig_139 <= '0';
      sig_140 <= '0';
      sig_141 <= '0';
      sig_142 <= '0';
      sig_143 <= '0';
      sig_144 <= '0';
      sig_145 <= '0';
      sig_146 <= '0';
      sig_147 <= '0';
      sig_148 <= '0';
      sig_149 <= '0';
      sig_150 <= '0';
      sig_151 <= '0';
      sig_152 <= '0';
      sig_153 <= '0';
      sig_154 <= '0';
      sig_155 <= '0';
      sig_156 <= '0';
      sig_157 <= '0';
      sig_158 <= '0';
      sig_159 <= '0';
      sig_160 <= '0';
      sig_161 <= '0';
      sig_162 <= '0';
      sig_163 <= '0';
      sig_164 <= '0';
      sig_165 <= '0';
      sig_166 <= '0';
      sig_167 <= '0';
      sig_168 <= '0';
      sig_169 <= '0';
      sig_170 <= '0';
      sig_171 <= '0';
      if (reg_start = '1') then
         sig_78 <= '1';
      else
         sig_78 <= '0';
      end if;
      if (reg_start = '1') then
         sig_79 <= '1';
      else
         sig_79 <= '0';
      end if;
      if (reg_next = '1') then
         sig_80 <= '1';
      else
         sig_80 <= '0';
      end if;
      if (reg_start = '1') then
         sig_81 <= '1';
      else
         sig_81 <= '0';
      end if;
      if (reg_next = '1') then
         sig_82 <= '1';
      else
         sig_82 <= '0';
      end if;
      if (reg_start = '1') then
         sig_83 <= '1';
      else
         sig_83 <= '0';
      end if;
      if (reg_next = '1') then
         sig_84 <= '1';
      else
         sig_84 <= '0';
      end if;
      if (reg_start = '1') then
         sig_85 <= '1';
      else
         sig_85 <= '0';
      end if;
      if (unsigned(reg_counter_misc) = 3) then
         sig_86 <= '1';
      else
         sig_86 <= '0';
      end if;
      if (unsigned(reg_counter_miller) = 0) then
         sig_87 <= '1';
      else
         sig_87 <= '0';
      end if;
      if (reg_add = '1') then
         sig_88 <= '1';
      else
         sig_88 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_89 <= '1';
      else
         sig_89 <= '0';
      end if;
      if (unsigned(reg_counter_miller) = 82) then
         sig_90 <= '1';
      else
         sig_90 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_91 <= '1';
      else
         sig_91 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_92 <= '1';
      else
         sig_92 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_93 <= '1';
      else
         sig_93 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_94 <= '1';
      else
         sig_94 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_95 <= '1';
      else
         sig_95 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_96 <= '1';
      else
         sig_96 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_97 <= '1';
      else
         sig_97 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_98 <= '1';
      else
         sig_98 <= '0';
      end if;
      if (unsigned(reg_counter_misc) = 5) then
         sig_99 <= '1';
      else
         sig_99 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_100 <= '1';
      else
         sig_100 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_101 <= '1';
      else
         sig_101 <= '0';
      end if;
      if (unsigned(reg_counter_misc) = 10) then
         sig_102 <= '1';
      else
         sig_102 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_103 <= '1';
      else
         sig_103 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_104 <= '1';
      else
         sig_104 <= '0';
      end if;
      if (unsigned(reg_counter_misc) = 20) then
         sig_105 <= '1';
      else
         sig_105 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_106 <= '1';
      else
         sig_106 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_107 <= '1';
      else
         sig_107 <= '0';
      end if;
      if (unsigned(reg_counter_misc) = 40) then
         sig_108 <= '1';
      else
         sig_108 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_109 <= '1';
      else
         sig_109 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_110 <= '1';
      else
         sig_110 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_111 <= '1';
      else
         sig_111 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_112 <= '1';
      else
         sig_112 <= '0';
      end if;
      if (unsigned(reg_counter_misc) = 81) then
         sig_113 <= '1';
      else
         sig_113 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_114 <= '1';
      else
         sig_114 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_115 <= '1';
      else
         sig_115 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_116 <= '1';
      else
         sig_116 <= '0';
      end if;
      if (unsigned(reg_counter_miller) = 0) then
         sig_117 <= '1';
      else
         sig_117 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_118 <= '1';
      else
         sig_118 <= '0';
      end if;
      if (reg_add = '0') then
         sig_119 <= '1';
      else
         sig_119 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_120 <= '1';
      else
         sig_120 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_121 <= '1';
      else
         sig_121 <= '0';
      end if;
      if (reg_add = '0') then
         sig_122 <= '1';
      else
         sig_122 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_123 <= '1';
      else
         sig_123 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_124 <= '1';
      else
         sig_124 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_125 <= '1';
      else
         sig_125 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_126 <= '1';
      else
         sig_126 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_127 <= '1';
      else
         sig_127 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_128 <= '1';
      else
         sig_128 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_129 <= '1';
      else
         sig_129 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_130 <= '1';
      else
         sig_130 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_131 <= '1';
      else
         sig_131 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_132 <= '1';
      else
         sig_132 <= '0';
      end if;
      if (unsigned(reg_counter_miller) = 82) then
         sig_133 <= '1';
      else
         sig_133 <= '0';
      end if;
      if (reg_add = '0') then
         sig_134 <= '1';
      else
         sig_134 <= '0';
      end if;
      sig_135 <= sig_133 and sig_134;
      if (reg_MALU_ready = '0') then
         sig_136 <= '1';
      else
         sig_136 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_137 <= '1';
      else
         sig_137 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_138 <= '1';
      else
         sig_138 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_139 <= '1';
      else
         sig_139 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_140 <= '1';
      else
         sig_140 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_141 <= '1';
      else
         sig_141 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_142 <= '1';
      else
         sig_142 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_143 <= '1';
      else
         sig_143 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_144 <= '1';
      else
         sig_144 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_145 <= '1';
      else
         sig_145 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_146 <= '1';
      else
         sig_146 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_147 <= '1';
      else
         sig_147 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_148 <= '1';
      else
         sig_148 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_149 <= '1';
      else
         sig_149 <= '0';
      end if;
      if (unsigned(reg_counter_misc) = 82) then
         sig_150 <= '1';
      else
         sig_150 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_151 <= '1';
      else
         sig_151 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_152 <= '1';
      else
         sig_152 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_153 <= '1';
      else
         sig_153 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_154 <= '1';
      else
         sig_154 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_155 <= '1';
      else
         sig_155 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_156 <= '1';
      else
         sig_156 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_157 <= '1';
      else
         sig_157 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_158 <= '1';
      else
         sig_158 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_159 <= '1';
      else
         sig_159 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_160 <= '1';
      else
         sig_160 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_161 <= '1';
      else
         sig_161 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_162 <= '1';
      else
         sig_162 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_163 <= '1';
      else
         sig_163 <= '0';
      end if;
      if (unsigned(reg_counter_misc) = 3) then
         sig_164 <= '1';
      else
         sig_164 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_165 <= '1';
      else
         sig_165 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_166 <= '1';
      else
         sig_166 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_167 <= '1';
      else
         sig_167 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_168 <= '1';
      else
         sig_168 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_169 <= '1';
      else
         sig_169 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_170 <= '1';
      else
         sig_170 <= '0';
      end if;
      if (reg_MALU_ready = '0') then
         sig_171 <= '1';
      else
         sig_171 <= '0';
      end if;
      cmd <= do_alwaysset_not_readyMALU_idleidle_ToMALUupdate_Xv_from_Inputidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
      case STATE is
         when init1 => 
            if (sig_78 = '1') then
                    cmd <= do_alwaysset_not_readyMALU_idleidle_ToMALUupdate_Xv_from_Inputidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleidle_regs;
            end if;
         when init2 => 
            if (sig_79 = '1') then
                    cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Inputidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
               if (sig_80 = '1') then
                       cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Inputupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
               else
                       cmd <= do_alwaysMALU_idleidle_regs;
               end if;
            end if;
         when init3 => 
            if (sig_81 = '1') then
                    cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Inputidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
               if (sig_82 = '1') then
                       cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Inputupdate_Yv_from_Xvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
               else
                       cmd <= do_alwaysMALU_idleidle_regs;
               end if;
            end if;
         when init4 => 
            if (sig_83 = '1') then
                    cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Inputidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
               if (sig_84 = '1') then
                       cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_Inputupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
               else
                       cmd <= do_alwaysMALU_idleidle_regs;
               end if;
            end if;
         when start => 
                 cmd <= do_alwaysMALU_addidle_regs;
         when distort1 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when distort2 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when distort3 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when distort4 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when distort5 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when distort6 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when distort7 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when distort8 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when miller_init1 => 
                 cmd <= do_alwaysMALU_idleunset_addreset_Freset_counter_milleridle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when miller_init2 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when startloop1 => 
            if (sig_87 = '1') then
                    cmd <= do_alwaysMALU_idleidle_regs;
            else
               if (sig_88 = '1') then
                       cmd <= do_alwaysMALU_idleidle_regs;
               else
                       cmd <= do_alwaysMALU_idleidle_regsdec_counter_miller;
               end if;
            end if;
         when ready1 => 
                 cmd <= do_alwaysset_readyreset_counter_miscMALU_idleidle_regs;
         when ready2 => 
            if (sig_85 = '1') then
                    cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Inputidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
               if (sig_86 = '1') then
                       cmd <= do_alwaysready_regsMALU_idle;
               else
                       cmd <= do_alwaysready_regsMALU_idle;
               end if;
            end if;
         when dlambda1 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when dlambda2 => 
                 cmd <= do_alwaysMALU_mult_plus_oneidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_Xv;
         when dlambda3 => 
            if (sig_89 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaupdate_Gb_from_Faupdate_Fa_from_Fbupdate_Fb_from_Fcupdate_Fc_from_Fdidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
            end if;
         when dlambda4 => 
            if (sig_90 = '1') then
                    cmd <= do_alwaysMALU_idleidle_regsset_add;
            else
                    cmd <= do_alwaysMALU_idleidle_regs;
            end if;
         when s => 
         when alambda1 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when alambda2 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when alambda3 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when alambda4 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaupdate_Gb_from_Faupdate_Fa_from_Fbupdate_Fb_from_Fcupdate_Fc_from_Fdidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when alambda5 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBidle_TmpB;
         when alambda6 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAidle_TmpAidle_TmpB;
         when alambda7 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when alambda8 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when alambda9 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when alambda10 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when alambda11 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when alambda12 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_Fdupdate_TmpB_from_Xv;
         when alambda13 => 
            if (sig_91 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
            end if;
         when alambda14 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when alambda15 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when alambda16 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when alambda17 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv1 => 
                 cmd <= do_alwaysreset_counter_miscMALU_idleupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when inv2 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBidle_TmpB;
         when inv3 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv4 => 
            if (sig_92 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv5 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv6 => 
            if (sig_93 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv7 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv8 => 
            if (sig_94 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv9 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when inv10 => 
            if (sig_95 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv11 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv12 => 
            if (sig_96 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv13 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA;
         when inv14 => 
            if (sig_97 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv15 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv16 => 
            if (sig_98 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv17 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv18 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when inv19 => 
            if (sig_99 = '1') then
                    cmd <= do_alwaysMALU_idleidle_regsreset_counter_misc;
            else
                    cmd <= do_alwaysinc_counter_miscMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv20 => 
            if (sig_100 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv21 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv22 => 
            if (sig_101 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv23 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv24 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when inv25 => 
            if (sig_102 = '1') then
                    cmd <= do_alwaysMALU_idleidle_regsreset_counter_misc;
            else
                    cmd <= do_alwaysinc_counter_miscMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv26 => 
            if (sig_103 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv27 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv28 => 
            if (sig_104 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv29 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv30 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when inv31 => 
            if (sig_105 = '1') then
                    cmd <= do_alwaysMALU_idleidle_regsreset_counter_misc;
            else
                    cmd <= do_alwaysinc_counter_miscMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv32 => 
            if (sig_106 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv33 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv34 => 
            if (sig_107 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv35 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv36 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when inv37 => 
            if (sig_108 = '1') then
                    cmd <= do_alwaysMALU_idleidle_regsreset_counter_misc;
            else
                    cmd <= do_alwaysinc_counter_miscMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv38 => 
            if (sig_109 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv39 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv40 => 
            if (sig_110 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv41 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA;
         when inv42 => 
            if (sig_111 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv43 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv44 => 
            if (sig_112 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv45 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv46 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when inv47 => 
            if (sig_113 = '1') then
                    cmd <= do_alwaysMALU_idleidle_regsreset_counter_misc;
            else
                    cmd <= do_alwaysinc_counter_miscMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv48 => 
            if (sig_114 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv49 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv50 => 
            if (sig_115 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv51 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv52 => 
            if (sig_116 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when inv53 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when inv54 => 
            if (sig_117 = '1') then
                    cmd <= do_alwaysMALU_idleidle_regs;
            else
                    cmd <= do_alwaysMALU_idleidle_regs;
            end if;
         when coord1 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when coord2 => 
            if (sig_118 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when coord3 => 
            if (sig_119 = '1') then
                    cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv;
            else
                    cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv;
            end if;
         when coord4 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when coord5 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when coord6 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when coord7 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when coord8 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when coord9 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when coord10 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv;
         when coord11 => 
            if (sig_120 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
            end if;
         when coord12 => 
                 cmd <= do_alwaysMALU_add_plus_oneidle_ToMALUupdate_Xv_from_TmpBidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when coord13 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when coord14 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when coord15 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when coord16 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when coord17 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when coord18 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when coord19 => 
            if (sig_121 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
            end if;
         when coord20 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when coord21 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when coord22 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when coord23 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when coord24 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when coord25 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when coord26 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when coord27 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Gbupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA;
         when coord28 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when coord29 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when coord30 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when coord31 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when coord32 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xvupdate_Xp_from_Yvidle_Ypupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA;
         when coord33 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdidle_TmpB;
         when coord34 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaupdate_Gb_from_Gaidle_Faidle_Fbupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA;
         when coord35 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when updatef1 => 
            if (sig_122 = '1') then
                    cmd <= do_alwaysMALU_idleidle_regs;
            else
                    cmd <= do_alwaysMALU_idleidle_regs;
            end if;
         when fsqrt1 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fsqrt2 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv;
         when fsqrt3 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fsqrt4 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fsqrt5 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when fsqrt6 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fsqrt7 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when fsqrt8 => 
            if (sig_123 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when fsqrt9 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when fsqrt10 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fsqrt11 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fsqrt12 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fsqrt13 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when fsqrt14 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when fsqrt15 => 
            if (sig_124 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when fsqrt16 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fsqrt17 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fsqrt18 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when fsqrt19 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fsqrt20 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fsqrt21 => 
                 cmd <= do_alwaysMALU_multupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when fsqrt22 => 
            if (sig_125 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
            end if;
         when fsqrt23 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when fsqrt24 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fsqrt25 => 
                 cmd <= do_alwaysMALU_multupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when fsqrt26 => 
            if (sig_126 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when fsqrt27 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fsqrt28 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fsqrt29 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB;
         when fsqrt30 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when fsqrt31 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fsqrt32 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fg1 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB;
         when fg2 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv;
         when fg3 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fg4 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fg5 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fg6 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when fg7 => 
            if (sig_127 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when fg8 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB;
         when fg9 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when fg10 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv;
         when fg11 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Fcupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv;
         when fg12 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when fg13 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fg14 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when fg15 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fg16 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when fg17 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fg18 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when fg19 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fg20 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fg21 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when fg22 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv;
         when fg23 => 
            if (sig_128 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
            end if;
         when fg24 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when fg25 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fg26 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fg27 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fg28 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when fg29 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fg30 => 
            if (sig_129 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
            end if;
         when fg31 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv;
         when fg32 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fg33 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when fg34 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fg35 => 
            if (sig_130 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
            end if;
         when fg36 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv;
         when fg37 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fg38 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when fg39 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fg40 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fg41 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv;
         when fg42 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fg43 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fg44 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fg45 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when fg46 => 
            if (sig_131 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
            end if;
         when fg47 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when fg48 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fg49 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA;
         when fg50 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when fg51 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when fg52 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_Fdupdate_TmpB_from_TmpA;
         when fg53 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fg54 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when fg55 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when fg56 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA;
         when fg57 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when fg58 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fg59 => 
            if (sig_132 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when fg60 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when fg61 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when fg62 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when fg63 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaupdate_Ga_from_Gbupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_Xv;
         when fg64 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_TmpBidle_TmpB;
         when fg65 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaupdate_Yfa_from_Gaupdate_Ga_from_Gbidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_TmpAidle_TmpAidle_TmpB;
         when fg66 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaupdate_Yfa_from_Gaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB;
         when fg67 => 
            if (sig_135 = '1') then
                    cmd <= do_alwaysMALU_idleidle_regsset_add;
            else
                    cmd <= unset_adddo_alwaysMALU_idleidle_regs;
            end if;
         when finalexp1 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdidle_TmpB;
         when finalexp2 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA;
         when finalexp3 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA;
         when finalexp4 => 
                 cmd <= do_alwaysMALU_multupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp5 => 
            if (sig_136 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when finalexp6 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp7 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when finalexp8 => 
                 cmd <= do_alwaysMALU_multupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when finalexp9 => 
            if (sig_137 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when finalexp10 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when finalexp11 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when finalexp12 => 
                 cmd <= do_alwaysMALU_multupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when finalexp13 => 
            if (sig_138 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when finalexp14 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp15 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when finalexp16 => 
                 cmd <= do_alwaysMALU_multupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp17 => 
            if (sig_139 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when finalexp18 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when finalexp19 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when finalexp20 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when finalexp21 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA;
         when finalexp22 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp23 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp24 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when finalexp25 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp26 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp27 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp28 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp29 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv;
         when finalexp30 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when finalexp31 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv;
         when finalexp32 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB;
         when finalexp33 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBidle_TmpB;
         when finalexp34 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp35 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when finalexp36 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp37 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp38 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Fcupdate_Fc_from_Fdupdate_Fd_from_TmpAidle_TmpAupdate_TmpB_from_Xv;
         when finalexp39 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBidle_TmpB;
         when finalexp40 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when finalexp41 => 
            if (sig_140 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when finalexp42 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp43 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp44 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp45 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when finalexp46 => 
            if (sig_141 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when finalexp47 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp48 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when finalexp49 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when finalexp50 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA;
         when finalexp51 => 
            if (sig_142 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when finalexp52 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp53 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp54 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp55 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp56 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Ypidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when finalexp57 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp58 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp59 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp60 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp61 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp62 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp63 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpupdate_Yp_from_Xpupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp64 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdidle_TmpB;
         when finalexp65 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAupdate_TmpB_from_TmpA;
         when finalexp66 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdidle_TmpB;
         when finalexp67 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA;
         when finalexp68 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_Fdupdate_TmpB_from_TmpA;
         when finalexp69 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp70 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp71 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when finalexp72 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when finalexp73 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp74 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp75 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Ypupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAidle_TmpAidle_TmpB;
         when finalexp76 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaupdate_Yfa_from_Xfaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when finalexp77 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaupdate_Ga_from_Yfaupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp78 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaupdate_Ga_from_Gbupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when finalexp79 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaupdate_Gb_from_Gaupdate_Fa_from_Gbupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcidle_TmpAidle_TmpB;
         when finalexp80 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Gbupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdidle_TmpB;
         when f4mpow1 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaupdate_Gb_from_Faupdate_Fa_from_Gbidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow2 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaupdate_Ga_from_Gbupdate_Gb_from_Gaupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow3 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaupdate_Yfa_from_Gaupdate_Ga_from_Yfaupdate_Gb_from_Faupdate_Fa_from_Gbidle_Fbupdate_Fc_from_Fbidle_Fdidle_TmpAidle_TmpB;
         when f4mpow4 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaupdate_Ga_from_Gbupdate_Gb_from_Gaupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcupdate_Fd_from_Fcidle_TmpAidle_TmpB;
         when f4mpow5 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faupdate_Fc_from_Fbidle_Fdidle_TmpAidle_TmpB;
         when f4mpow6 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaupdate_Gb_from_Faupdate_Fa_from_Gbidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow7 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaupdate_Ga_from_Gbupdate_Gb_from_Gaupdate_Fa_from_Fbupdate_Fb_from_Faidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow8 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaupdate_Gb_from_Faupdate_Fa_from_Gbidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow9 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow10 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xfaidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow11 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Ypidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow12 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow13 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow14 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow15 => 
            if (sig_143 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when f4mpow16 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaupdate_Ga_from_Gbupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow17 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow18 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaupdate_Ga_from_Gbupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when f4mpow19 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xfaidle_Xfaupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow20 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBidle_TmpB;
         when f4mpow21 => 
            if (sig_144 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
            end if;
         when f4mpow22 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xfaidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow23 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow24 => 
            if (sig_145 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when f4mpow25 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow26 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow27 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow28 => 
            if (sig_146 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when f4mpow29 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow30 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow31 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow32 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow33 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow34 => 
            if (sig_147 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when f4mpow35 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow36 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when f4mpow37 => 
            if (sig_148 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when f4mpow38 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow39 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow40 => 
            if (sig_149 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when f4mpow41 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow42 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow43 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when f4mpow44 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow45 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow46 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow47 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when f4mpow48 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow49 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow50 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow51 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow52 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow53 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA;
         when f4mpow54 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow55 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow56 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaupdate_Yfa_from_Xfaupdate_Ga_from_Yfaupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow57 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow58 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaupdate_Yfa_from_Gaupdate_Ga_from_Yfaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow59 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaupdate_Ga_from_Gbupdate_Gb_from_Gaidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow60 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mpow61 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdidle_TmpB;
         when f4mpow62 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA;
         when f4mpow47fix => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt1 => 
                 cmd <= do_alwaysMALU_idleidle_regsreset_counter_misc;
         when f4msqrt2 => 
            if (sig_150 = '1') then
                    cmd <= do_alwaysMALU_idleidle_regsreset_counter_misc;
            else
                    cmd <= do_alwaysinc_counter_miscMALU_idleidle_regs;
            end if;
         when f4msqrt3 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA;
         when f4msqrt4 => 
                 cmd <= do_alwaysMALU_multupdate_ToMALU_from_Xvidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt5 => 
            if (sig_151 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_Fdupdate_TmpB_from_TmpA;
            end if;
         when f4msqrt6 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt7 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt8 => 
            if (sig_152 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA;
            end if;
         when f4msqrt9 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt10 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt11 => 
            if (sig_153 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when f4msqrt12 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt13 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt14 => 
            if (sig_154 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when f4msqrt15 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt16 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Ypidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt17 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt18 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt19 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt20 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt21 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt22 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt23 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt24 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt25 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4msqrt26 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_Xv;
         when f4msqrt27 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv;
         when f4msqrt28 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_Xv;
         when f4msqrt29 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f4msqrt30 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when f4msqrt31 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f4msqrt32 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when f4msqrt27fix => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_Xv;
         when f4mmult1 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Yfaupdate_Yfa_from_Gaupdate_Ga_from_Gbidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f4mmult2 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_TmpBupdate_Yv_from_Xvupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaupdate_Yfa_from_Gaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when f4mmult3 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f4mmult4 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult5 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult6 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult7 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult8 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult9 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Ypupdate_Yp_from_Xpupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult10 => 
            if (sig_155 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_TmpBidle_TmpB;
            end if;
         when f4mmult11 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when f4mmult12 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult13 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when f4mmult14 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult15 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypupdate_Xfa_from_Yfaupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBidle_TmpB;
         when f4mmult16 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv;
         when f4mmult17 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f4mmult18 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv;
         when f4mmult19 => 
            if (sig_156 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
            end if;
         when f4mmult20 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when f4mmult21 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult22 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbidle_Fdidle_TmpAidle_TmpB;
         when f4mmult23 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB;
         when f4mmult24 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv;
         when f4mmult25 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f4mmult26 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv;
         when f4mmult27 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f4mmult28 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Fcupdate_Fc_from_Fdupdate_Fd_from_TmpAupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f4mmult29 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaupdate_Gb_from_Faupdate_Fa_from_Fbupdate_Fb_from_Faupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAupdate_TmpB_from_Xv;
         when f4mmult30 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f4mmult31 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAupdate_TmpB_from_Xv;
         when f4mmult32 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f4mmult33 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when f4mmult34 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f4mmult35 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAupdate_TmpB_from_Xv;
         when f4mmult36 => 
            if (sig_157 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
            end if;
         when f4mmult37 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv;
         when f4mmult38 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f4mmult39 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when f4mmult40 => 
            if (sig_158 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
            end if;
         when f4mmult41 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when f4mmult42 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when f4mmult43 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f4mmult44 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when f4mmult45 => 
            if (sig_159 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Faupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAupdate_TmpB_from_TmpA;
            end if;
         when f4mmult46 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Fcupdate_Fc_from_Fbidle_Fdupdate_TmpA_from_Fdidle_TmpB;
         when f4mmult47 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_Fcidle_TmpAidle_TmpB;
         when f4mmult48 => 
            if (sig_160 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
            end if;
         when f4mmult49 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult50 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when f4mmult51 => 
            if (sig_161 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
            end if;
         when f4mmult52 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f4mmult53 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when f4mmult54 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult55 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult56 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when f4mmult57 => 
            if (sig_162 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
            end if;
         when f4mmult58 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult59 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Faupdate_Fc_from_Fbidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when f4mmult60 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbupdate_Fc_from_Fdupdate_Fd_from_Fcidle_TmpAidle_TmpB;
         when f4mmult61 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbupdate_Fa_from_Fbupdate_Fb_from_Fcupdate_Fc_from_Fbupdate_Fd_from_TmpAupdate_TmpA_from_Fdidle_TmpB;
         when f4mmult62 => 
            if (sig_163 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_Fdupdate_TmpB_from_TmpA;
            end if;
         when f4mmult63 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult64 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f4mmult65 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult66 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcidle_TmpAidle_TmpB;
         when f4mmult67 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv;
         when f4mmult68 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpupdate_Yp_from_Xfaupdate_Xfa_from_Ypupdate_Yfa_from_Xfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f4mmult69 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult70 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when f4mmult71 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult72 => 
         when f4mmult73 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult74 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult75 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult76 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult77 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult78 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult79 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult80 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult81 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult82 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA;
         when f4mmult83 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcupdate_Fd_from_TmpAupdate_TmpA_from_Fdupdate_TmpB_from_Xv;
         when f4mmult84 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f4mmult85 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_Fdupdate_TmpB_from_TmpA;
         when f4mmult86 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f4mmult87 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Ypidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult88 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult89 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult90 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult91 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA;
         when f4mmult92 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult93 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult94 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult95 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmult96 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmfix1 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmfix2 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmfix3 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvupdate_Yp_from_Xfaupdate_Xfa_from_Ypidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmfix4 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f4mmfix5 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xfaupdate_Xfa_from_Yfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2mmult1 => 
                 cmd <= do_alwaysMALU_idleidle_regsreset_counter_misc;
         when f2mmult2 => 
            if (sig_164 = '1') then
                    cmd <= do_alwaysMALU_idleidle_regsreset_counter_misc;
            else
                    cmd <= do_alwaysinc_counter_miscMALU_idleidle_regs;
            end if;
         when f2mmult3 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f2mmult4 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f2mmult5 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2mmult6 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2mmult7 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2mmult8 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2mmult9 => 
            if (sig_165 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when f2mmult10 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2mmult11 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xpupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when f2mmult12 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2mmult13 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdupdate_TmpA_from_TmpBupdate_TmpB_from_TmpA;
         when f2mmult14 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2mmult15 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when f2mmult16 => 
            if (sig_166 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_Yvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when f2mmult17 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2mmult18 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when f2mmult19 => 
            if (sig_167 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_TmpA;
            end if;
         when f2mmult20 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2mmult21 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2mmult22 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2mmult23 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_TmpBupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2mmult24 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2mmult25 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2mmult26 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvupdate_Xp_from_Ypupdate_Yp_from_Xpidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2mmult27 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xpupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2mmult28 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvupdate_Yv_from_Xvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaupdate_Gb_from_Gaupdate_Fa_from_Gbupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA;
         when f2mmult29 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUidle_Xvidle_Yvupdate_Xp_from_Yvupdate_Yp_from_Xpupdate_Xfa_from_Ypupdate_Yfa_from_Xfaupdate_Ga_from_Yfaupdate_Gb_from_Gaupdate_Fa_from_Gbupdate_Fb_from_Faupdate_Fc_from_Fbupdate_Fd_from_Fcupdate_TmpA_from_Fdupdate_TmpB_from_TmpA;
         when f2minv1 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2minv2 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2minv3 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2minv4 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2minv5 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when f2minv6 => 
            if (sig_168 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when f2minv7 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvupdate_Xp_from_Yvidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2minv8 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2minv9 => 
                 cmd <= do_alwaysMALU_multupdate_ToMALU_from_Xvupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2minv10 => 
            if (sig_169 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when f2minv11 => 
                 cmd <= do_alwaysMALU_addidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2minv12 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2minv13 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2minv14 => 
                 cmd <= do_alwaysMALU_multupdate_ToMALU_from_Xvupdate_Xv_from_Yvupdate_Yv_from_Xpidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAupdate_TmpB_from_Xv;
         when f2minv15 => 
            if (sig_170 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUupdate_Xv_from_TmpBidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when f2minv16 => 
                 cmd <= do_alwaysMALU_idleupdate_ToMALU_from_Xvupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2minv17 => 
                 cmd <= do_alwaysMALU_multidle_ToMALUupdate_Xv_from_Yvupdate_Yv_from_Xvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when f2minv18 => 
            if (sig_171 = '1') then
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_ToMALUShiftidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            else
                    cmd <= do_alwaysMALU_idleupdate_ToMALU_from_MALUidle_Xvidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
            end if;
         when f2minv19 => 
                 cmd <= do_alwaysMALU_idleidle_ToMALUupdate_Xv_from_ToMALUidle_Yvidle_Xpidle_Ypidle_Xfaidle_Yfaidle_Gaidle_Gbidle_Faidle_Fbidle_Fcidle_Fdidle_TmpAidle_TmpB;
         when others=>
         end case;
   end process fsmCMB;

	CLK_Xv <= CLK and sig_en_Xv;
	CLK_Yv <= CLK and sig_en_Yv;
	CLK_Xp <= CLK and sig_en_Xp;
	CLK_Yp <= CLK and sig_en_Yp;
	CLK_Xfa <= CLK and sig_en_Xfa;
	CLK_Yfa <= CLK and sig_en_Yfa;
	CLK_Ga <= CLK and sig_en_Ga;
	CLK_Gb <= CLK and sig_en_Gb;
	CLK_Fa <= CLK and sig_en_Fa;
	CLK_Fb <= CLK and sig_en_Fb;
	CLK_Fc <= CLK and sig_en_Fc;
	CLK_Fd <= CLK and sig_en_Fd;
	CLK_TmpA <= CLK and sig_en_TmpA;
	CLK_TmpB <= CLK and sig_en_TmpB;
	CLK_ToMALU <= CLK and sig_en_ToMALU;
end RTL;
